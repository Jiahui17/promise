module iterative_division(
  input [7:0] dividend,
  input  dividend_valid,
  input [7:0] divisor,
  input  divisor_valid,
  input  start_valid,
  input  clk,
  input  rst,
  input  out0_ready,
  input  end_ready,
  output  dividend_ready,
  output  divisor_ready,
  output  start_ready,
  output [7:0] out0,
  output  out0_valid,
  output  end_valid
);
  wire  fork0_outs_0_valid;
  wire  fork0_outs_0_ready;
  wire  fork0_outs_1_valid;
  wire  fork0_outs_1_ready;
  wire  fork0_outs_2_valid;
  wire  fork0_outs_2_ready;
  wire [7:0] fork1_outs_0;
  wire  fork1_outs_0_valid;
  wire  fork1_outs_0_ready;
  wire [7:0] fork1_outs_1;
  wire  fork1_outs_1_valid;
  wire  fork1_outs_1_ready;
  wire [7:0] fork1_outs_2;
  wire  fork1_outs_2_valid;
  wire  fork1_outs_2_ready;
  wire  source0_outs_valid;
  wire  source0_outs_ready;
  wire [0:0] constant1_outs;
  wire  constant1_outs_valid;
  wire  constant1_outs_ready;
  wire [0:0] fork2_outs_0;
  wire  fork2_outs_0_valid;
  wire  fork2_outs_0_ready;
  wire [0:0] fork2_outs_1;
  wire  fork2_outs_1_valid;
  wire  fork2_outs_1_ready;
  wire [7:0] extsi15_outs;
  wire  extsi15_outs_valid;
  wire  extsi15_outs_ready;
  wire [7:0] extsi16_outs;
  wire  extsi16_outs_valid;
  wire  extsi16_outs_ready;
  wire [0:0] constant2_outs;
  wire  constant2_outs_valid;
  wire  constant2_outs_ready;
  wire [0:0] cmpi0_result;
  wire  cmpi0_result_valid;
  wire  cmpi0_result_ready;
  wire [0:0] cmpi1_result;
  wire  cmpi1_result_valid;
  wire  cmpi1_result_ready;
  wire [0:0] fork3_outs_0;
  wire  fork3_outs_0_valid;
  wire  fork3_outs_0_ready;
  wire [0:0] fork3_outs_1;
  wire  fork3_outs_1_valid;
  wire  fork3_outs_1_ready;
  wire [0:0] fork3_outs_2;
  wire  fork3_outs_2_valid;
  wire  fork3_outs_2_ready;
  wire [0:0] fork3_outs_3;
  wire  fork3_outs_3_valid;
  wire  fork3_outs_3_ready;
  wire [0:0] fork3_outs_4;
  wire  fork3_outs_4_valid;
  wire  fork3_outs_4_ready;
  wire [7:0] cond_br3_trueOut;
  wire  cond_br3_trueOut_valid;
  wire  cond_br3_trueOut_ready;
  wire [7:0] cond_br3_falseOut;
  wire  cond_br3_falseOut_valid;
  wire  cond_br3_falseOut_ready;
  wire [7:0] cond_br4_trueOut;
  wire  cond_br4_trueOut_valid;
  wire  cond_br4_trueOut_ready;
  wire [7:0] cond_br4_falseOut;
  wire  cond_br4_falseOut_valid;
  wire  cond_br4_falseOut_ready;
  wire  cond_br5_trueOut_valid;
  wire  cond_br5_trueOut_ready;
  wire  cond_br5_falseOut_valid;
  wire  cond_br5_falseOut_ready;
  wire [0:0] cond_br6_trueOut;
  wire  cond_br6_trueOut_valid;
  wire  cond_br6_trueOut_ready;
  wire [0:0] cond_br6_falseOut;
  wire  cond_br6_falseOut_valid;
  wire  cond_br6_falseOut_ready;
  wire [0:0] cond_br7_trueOut;
  wire  cond_br7_trueOut_valid;
  wire  cond_br7_trueOut_ready;
  wire [0:0] cond_br7_falseOut;
  wire  cond_br7_falseOut_valid;
  wire  cond_br7_falseOut_ready;
  wire [7:0] buffer0_outs;
  wire  buffer0_outs_valid;
  wire  buffer0_outs_ready;
  wire [7:0] buffer1_outs;
  wire  buffer1_outs_valid;
  wire  buffer1_outs_ready;
  wire [7:0] fork4_outs_0;
  wire  fork4_outs_0_valid;
  wire  fork4_outs_0_ready;
  wire [7:0] fork4_outs_1;
  wire  fork4_outs_1_valid;
  wire  fork4_outs_1_ready;
  wire [7:0] fork4_outs_2;
  wire  fork4_outs_2_valid;
  wire  fork4_outs_2_ready;
  wire [7:0] fork4_outs_3;
  wire  fork4_outs_3_valid;
  wire  fork4_outs_3_ready;
  wire [7:0] buffer2_outs;
  wire  buffer2_outs_valid;
  wire  buffer2_outs_ready;
  wire [7:0] buffer3_outs;
  wire  buffer3_outs_valid;
  wire  buffer3_outs_ready;
  wire [7:0] fork5_outs_0;
  wire  fork5_outs_0_valid;
  wire  fork5_outs_0_ready;
  wire [7:0] fork5_outs_1;
  wire  fork5_outs_1_valid;
  wire  fork5_outs_1_ready;
  wire [7:0] fork5_outs_2;
  wire  fork5_outs_2_valid;
  wire  fork5_outs_2_ready;
  wire [7:0] fork5_outs_3;
  wire  fork5_outs_3_valid;
  wire  fork5_outs_3_ready;
  wire  buffer4_outs_valid;
  wire  buffer4_outs_ready;
  wire  buffer5_outs_valid;
  wire  buffer5_outs_ready;
  wire  fork6_outs_0_valid;
  wire  fork6_outs_0_ready;
  wire  fork6_outs_1_valid;
  wire  fork6_outs_1_ready;
  wire  source1_outs_valid;
  wire  source1_outs_ready;
  wire [1:0] constant3_outs;
  wire  constant3_outs_valid;
  wire  constant3_outs_ready;
  wire [7:0] extsi17_outs;
  wire  extsi17_outs_valid;
  wire  extsi17_outs_ready;
  wire  source2_outs_valid;
  wire  source2_outs_ready;
  wire [31:0] constant7_outs;
  wire  constant7_outs_valid;
  wire  constant7_outs_ready;
  wire [7:0] trunci5_outs;
  wire  trunci5_outs_valid;
  wire  trunci5_outs_ready;
  wire [0:0] constant4_outs;
  wire  constant4_outs_valid;
  wire  constant4_outs_ready;
  wire  source3_outs_valid;
  wire  source3_outs_ready;
  wire [0:0] constant5_outs;
  wire  constant5_outs_valid;
  wire  constant5_outs_ready;
  wire [0:0] fork7_outs_0;
  wire  fork7_outs_0_valid;
  wire  fork7_outs_0_ready;
  wire [0:0] fork7_outs_1;
  wire  fork7_outs_1_valid;
  wire  fork7_outs_1_ready;
  wire [0:0] fork7_outs_2;
  wire  fork7_outs_2_valid;
  wire  fork7_outs_2_ready;
  wire [0:0] fork7_outs_3;
  wire  fork7_outs_3_valid;
  wire  fork7_outs_3_ready;
  wire [0:0] fork7_outs_4;
  wire  fork7_outs_4_valid;
  wire  fork7_outs_4_ready;
  wire [0:0] fork7_outs_5;
  wire  fork7_outs_5_valid;
  wire  fork7_outs_5_ready;
  wire [7:0] extsi18_outs;
  wire  extsi18_outs_valid;
  wire  extsi18_outs_ready;
  wire [7:0] extsi19_outs;
  wire  extsi19_outs_valid;
  wire  extsi19_outs_ready;
  wire [7:0] extsi20_outs;
  wire  extsi20_outs_valid;
  wire  extsi20_outs_ready;
  wire [7:0] extsi21_outs;
  wire  extsi21_outs_valid;
  wire  extsi21_outs_ready;
  wire [7:0] extsi22_outs;
  wire  extsi22_outs_valid;
  wire  extsi22_outs_ready;
  wire [7:0] extsi23_outs;
  wire  extsi23_outs_valid;
  wire  extsi23_outs_ready;
  wire [0:0] cmpi2_result;
  wire  cmpi2_result_valid;
  wire  cmpi2_result_ready;
  wire [0:0] cmpi3_result;
  wire  cmpi3_result_valid;
  wire  cmpi3_result_ready;
  wire [0:0] xori0_result;
  wire  xori0_result_valid;
  wire  xori0_result_ready;
  wire [7:0] select0_result;
  wire  select0_result_valid;
  wire  select0_result_ready;
  wire [0:0] cmpi4_result;
  wire  cmpi4_result_valid;
  wire  cmpi4_result_ready;
  wire [7:0] subi4_result;
  wire  subi4_result_valid;
  wire  subi4_result_ready;
  wire [7:0] select2_result;
  wire  select2_result_valid;
  wire  select2_result_ready;
  wire [0:0] cmpi5_result;
  wire  cmpi5_result_valid;
  wire  cmpi5_result_ready;
  wire [7:0] subi5_result;
  wire  subi5_result_valid;
  wire  subi5_result_ready;
  wire [7:0] select3_result;
  wire  select3_result_valid;
  wire  select3_result_ready;
  wire [7:0] extsi24_outs;
  wire  extsi24_outs_valid;
  wire  extsi24_outs_ready;
  wire [7:0] mux0_outs;
  wire  mux0_outs_valid;
  wire  mux0_outs_ready;
  wire [7:0] mux1_outs;
  wire  mux1_outs_valid;
  wire  mux1_outs_ready;
  wire [7:0] buffer8_outs;
  wire  buffer8_outs_valid;
  wire  buffer8_outs_ready;
  wire [7:0] buffer9_outs;
  wire  buffer9_outs_valid;
  wire  buffer9_outs_ready;
  wire [7:0] fork8_outs_0;
  wire  fork8_outs_0_valid;
  wire  fork8_outs_0_ready;
  wire [7:0] fork8_outs_1;
  wire  fork8_outs_1_valid;
  wire  fork8_outs_1_ready;
  wire [7:0] mux2_outs;
  wire  mux2_outs_valid;
  wire  mux2_outs_ready;
  wire [7:0] mux3_outs;
  wire  mux3_outs_valid;
  wire  mux3_outs_ready;
  wire [7:0] buffer12_outs;
  wire  buffer12_outs_valid;
  wire  buffer12_outs_ready;
  wire [7:0] buffer13_outs;
  wire  buffer13_outs_valid;
  wire  buffer13_outs_ready;
  wire [7:0] fork9_outs_0;
  wire  fork9_outs_0_valid;
  wire  fork9_outs_0_ready;
  wire [7:0] fork9_outs_1;
  wire  fork9_outs_1_valid;
  wire  fork9_outs_1_ready;
  wire  control_merge1_outs_valid;
  wire  control_merge1_outs_ready;
  wire [0:0] control_merge1_index;
  wire  control_merge1_index_valid;
  wire  control_merge1_index_ready;
  wire [0:0] fork10_outs_0;
  wire  fork10_outs_0_valid;
  wire  fork10_outs_0_ready;
  wire [0:0] fork10_outs_1;
  wire  fork10_outs_1_valid;
  wire  fork10_outs_1_ready;
  wire [0:0] fork10_outs_2;
  wire  fork10_outs_2_valid;
  wire  fork10_outs_2_ready;
  wire [0:0] fork10_outs_3;
  wire  fork10_outs_3_valid;
  wire  fork10_outs_3_ready;
  wire [0:0] cmpi6_result;
  wire  cmpi6_result_valid;
  wire  cmpi6_result_ready;
  wire [0:0] fork11_outs_0;
  wire  fork11_outs_0_valid;
  wire  fork11_outs_0_ready;
  wire [0:0] fork11_outs_1;
  wire  fork11_outs_1_valid;
  wire  fork11_outs_1_ready;
  wire [0:0] fork11_outs_2;
  wire  fork11_outs_2_valid;
  wire  fork11_outs_2_ready;
  wire [0:0] fork11_outs_3;
  wire  fork11_outs_3_valid;
  wire  fork11_outs_3_ready;
  wire [0:0] fork11_outs_4;
  wire  fork11_outs_4_valid;
  wire  fork11_outs_4_ready;
  wire [7:0] buffer6_outs;
  wire  buffer6_outs_valid;
  wire  buffer6_outs_ready;
  wire [7:0] buffer7_outs;
  wire  buffer7_outs_valid;
  wire  buffer7_outs_ready;
  wire [7:0] cond_br8_trueOut;
  wire  cond_br8_trueOut_valid;
  wire  cond_br8_trueOut_ready;
  wire [7:0] cond_br8_falseOut;
  wire  cond_br8_falseOut_valid;
  wire  cond_br8_falseOut_ready;
  wire [7:0] cond_br9_trueOut;
  wire  cond_br9_trueOut_valid;
  wire  cond_br9_trueOut_ready;
  wire [7:0] cond_br9_falseOut;
  wire  cond_br9_falseOut_valid;
  wire  cond_br9_falseOut_ready;
  wire [7:0] buffer10_outs;
  wire  buffer10_outs_valid;
  wire  buffer10_outs_ready;
  wire [7:0] buffer11_outs;
  wire  buffer11_outs_valid;
  wire  buffer11_outs_ready;
  wire [7:0] cond_br10_trueOut;
  wire  cond_br10_trueOut_valid;
  wire  cond_br10_trueOut_ready;
  wire [7:0] cond_br10_falseOut;
  wire  cond_br10_falseOut_valid;
  wire  cond_br10_falseOut_ready;
  wire [7:0] cond_br11_trueOut;
  wire  cond_br11_trueOut_valid;
  wire  cond_br11_trueOut_ready;
  wire [7:0] cond_br11_falseOut;
  wire  cond_br11_falseOut_valid;
  wire  cond_br11_falseOut_ready;
  wire  buffer14_outs_valid;
  wire  buffer14_outs_ready;
  wire  buffer15_outs_valid;
  wire  buffer15_outs_ready;
  wire  cond_br12_trueOut_valid;
  wire  cond_br12_trueOut_ready;
  wire  cond_br12_falseOut_valid;
  wire  cond_br12_falseOut_ready;
  wire [7:0] buffer22_outs;
  wire  buffer22_outs_valid;
  wire  buffer22_outs_ready;
  wire [7:0] buffer23_outs;
  wire  buffer23_outs_valid;
  wire  buffer23_outs_ready;
  wire [7:0] fork12_outs_0;
  wire  fork12_outs_0_valid;
  wire  fork12_outs_0_ready;
  wire [7:0] fork12_outs_1;
  wire  fork12_outs_1_valid;
  wire  fork12_outs_1_ready;
  wire  source4_outs_valid;
  wire  source4_outs_ready;
  wire [1:0] constant14_outs;
  wire  constant14_outs_valid;
  wire  constant14_outs_ready;
  wire [7:0] extsi13_outs;
  wire  extsi13_outs_valid;
  wire  extsi13_outs_ready;
  wire [7:0] buffer18_outs;
  wire  buffer18_outs_valid;
  wire  buffer18_outs_ready;
  wire [7:0] buffer19_outs;
  wire  buffer19_outs_valid;
  wire  buffer19_outs_ready;
  wire [7:0] subi2_result;
  wire  subi2_result_valid;
  wire  subi2_result_ready;
  wire [7:0] buffer16_outs;
  wire  buffer16_outs_valid;
  wire  buffer16_outs_ready;
  wire [7:0] buffer17_outs;
  wire  buffer17_outs_valid;
  wire  buffer17_outs_ready;
  wire [7:0] addi0_result;
  wire  addi0_result_valid;
  wire  addi0_result_ready;
  wire [7:0] buffer20_outs;
  wire  buffer20_outs_valid;
  wire  buffer20_outs_ready;
  wire [7:0] buffer21_outs;
  wire  buffer21_outs_valid;
  wire  buffer21_outs_ready;
  wire  buffer24_outs_valid;
  wire  buffer24_outs_ready;
  wire  buffer25_outs_valid;
  wire  buffer25_outs_ready;
  wire  source5_outs_valid;
  wire  source5_outs_ready;
  wire [31:0] constant11_outs;
  wire  constant11_outs_valid;
  wire  constant11_outs_ready;
  wire [7:0] buffer26_outs;
  wire  buffer26_outs_valid;
  wire  buffer26_outs_ready;
  wire [7:0] buffer27_outs;
  wire  buffer27_outs_valid;
  wire  buffer27_outs_ready;
  wire [31:0] extsi5_outs;
  wire  extsi5_outs_valid;
  wire  extsi5_outs_ready;
  wire [0:0] cmpi7_result;
  wire  cmpi7_result_valid;
  wire  cmpi7_result_ready;
  wire [0:0] fork13_outs_0;
  wire  fork13_outs_0_valid;
  wire  fork13_outs_0_ready;
  wire [0:0] fork13_outs_1;
  wire  fork13_outs_1_valid;
  wire  fork13_outs_1_ready;
  wire [7:0] buffer28_outs;
  wire  buffer28_outs_valid;
  wire  buffer28_outs_ready;
  wire [7:0] buffer29_outs;
  wire  buffer29_outs_valid;
  wire  buffer29_outs_ready;
  wire [7:0] cond_br13_trueOut;
  wire  cond_br13_trueOut_valid;
  wire  cond_br13_trueOut_ready;
  wire [7:0] cond_br13_falseOut;
  wire  cond_br13_falseOut_valid;
  wire  cond_br13_falseOut_ready;
  wire  buffer30_outs_valid;
  wire  buffer30_outs_ready;
  wire  buffer31_outs_valid;
  wire  buffer31_outs_ready;
  wire  cond_br14_trueOut_valid;
  wire  cond_br14_trueOut_ready;
  wire  cond_br14_falseOut_valid;
  wire  cond_br14_falseOut_ready;
  wire  source6_outs_valid;
  wire  source6_outs_ready;
  wire [0:0] constant15_outs;
  wire  constant15_outs_valid;
  wire  constant15_outs_ready;
  wire [7:0] extsi25_outs;
  wire  extsi25_outs_valid;
  wire  extsi25_outs_ready;
  wire [7:0] buffer32_outs;
  wire  buffer32_outs_valid;
  wire  buffer32_outs_ready;
  wire [7:0] buffer33_outs;
  wire  buffer33_outs_valid;
  wire  buffer33_outs_ready;
  wire [7:0] subi3_result;
  wire  subi3_result_valid;
  wire  subi3_result_ready;
  wire  buffer34_outs_valid;
  wire  buffer34_outs_ready;
  wire  buffer35_outs_valid;
  wire  buffer35_outs_ready;
  wire [7:0] buffer36_outs;
  wire  buffer36_outs_valid;
  wire  buffer36_outs_ready;
  wire [7:0] buffer37_outs;
  wire  buffer37_outs_valid;
  wire  buffer37_outs_ready;
  wire  buffer38_outs_valid;
  wire  buffer38_outs_ready;
  wire  buffer39_outs_valid;
  wire  buffer39_outs_ready;
  wire [7:0] mux4_outs;
  wire  mux4_outs_valid;
  wire  mux4_outs_ready;
  wire  control_merge6_outs_valid;
  wire  control_merge6_outs_ready;
  wire [0:0] control_merge6_index;
  wire  control_merge6_index_valid;
  wire  control_merge6_index_ready;
  wire [7:0] buffer40_outs;
  wire  buffer40_outs_valid;
  wire  buffer40_outs_ready;
  wire [7:0] buffer41_outs;
  wire  buffer41_outs_valid;
  wire  buffer41_outs_ready;
  wire  buffer42_outs_valid;
  wire  buffer42_outs_ready;
  wire  buffer43_outs_valid;
  wire  buffer43_outs_ready;
  wire [0:0] buffer44_outs;
  wire  buffer44_outs_valid;
  wire  buffer44_outs_ready;
  wire [0:0] buffer45_outs;
  wire  buffer45_outs_valid;
  wire  buffer45_outs_ready;
  wire [7:0] extsi26_outs;
  wire  extsi26_outs_valid;
  wire  extsi26_outs_ready;
  wire  source7_outs_valid;
  wire  source7_outs_ready;
  wire [7:0] constant13_outs;
  wire  constant13_outs_valid;
  wire  constant13_outs_ready;
  wire [0:0] buffer46_outs;
  wire  buffer46_outs_valid;
  wire  buffer46_outs_ready;
  wire [0:0] buffer47_outs;
  wire  buffer47_outs_valid;
  wire  buffer47_outs_ready;
  wire [7:0] select1_result;
  wire  select1_result_valid;
  wire  select1_result_ready;
  wire  buffer48_outs_valid;
  wire  buffer48_outs_ready;
  wire  buffer49_outs_valid;
  wire  buffer49_outs_ready;
  wire [7:0] mux5_outs;
  wire  mux5_outs_valid;
  wire  mux5_outs_ready;
  wire  control_merge8_outs_valid;
  wire  control_merge8_outs_ready;
  wire [0:0] control_merge8_index;
  wire  control_merge8_index_valid;
  wire  control_merge8_index_ready;
  wire  buffer52_outs_valid;
  wire  buffer52_outs_ready;
  wire  buffer53_outs_valid;
  wire  buffer53_outs_ready;
  wire [7:0] buffer50_outs;
  wire  buffer50_outs_valid;
  wire  buffer50_outs_ready;
  wire [7:0] buffer51_outs;
  wire  buffer51_outs_valid;
  wire  buffer51_outs_ready;

  assign out0 = buffer51_outs;
  assign out0_valid = buffer51_outs_valid;
  assign buffer51_outs_ready = out0_ready;
  assign end_valid = fork0_outs_1_valid;
  assign fork0_outs_1_ready = end_ready;

  fork_dataless #(.SIZE(3)) fork0(
    .ins_valid (start_valid),
    .ins_ready (start_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork0_outs_2_valid, fork0_outs_1_valid, fork0_outs_0_valid}),
    .outs_ready ({fork0_outs_2_ready, fork0_outs_1_ready, fork0_outs_0_ready})
  );

  fork_type #(.SIZE(3), .DATA_TYPE(8)) fork1(
    .ins (divisor),
    .ins_valid (divisor_valid),
    .ins_ready (divisor_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork1_outs_2, fork1_outs_1, fork1_outs_0}),
    .outs_valid ({fork1_outs_2_valid, fork1_outs_1_valid, fork1_outs_0_valid}),
    .outs_ready ({fork1_outs_2_ready, fork1_outs_1_ready, fork1_outs_0_ready})
  );

  source source0(
    .clk (clk),
    .rst (rst),
    .outs_valid (source0_outs_valid),
    .outs_ready (source0_outs_ready)
  );

  handshake_constant_0 #(.DATA_WIDTH(1)) constant1(
    .ctrl_valid (source0_outs_valid),
    .ctrl_ready (source0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant1_outs),
    .outs_valid (constant1_outs_valid),
    .outs_ready (constant1_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(1)) fork2(
    .ins (constant1_outs),
    .ins_valid (constant1_outs_valid),
    .ins_ready (constant1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork2_outs_1, fork2_outs_0}),
    .outs_valid ({fork2_outs_1_valid, fork2_outs_0_valid}),
    .outs_ready ({fork2_outs_1_ready, fork2_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi15(
    .ins (fork2_outs_0),
    .ins_valid (fork2_outs_0_valid),
    .ins_ready (fork2_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi15_outs),
    .outs_valid (extsi15_outs_valid),
    .outs_ready (extsi15_outs_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi16(
    .ins (fork2_outs_1),
    .ins_valid (fork2_outs_1_valid),
    .ins_ready (fork2_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi16_outs),
    .outs_valid (extsi16_outs_valid),
    .outs_ready (extsi16_outs_ready)
  );

  handshake_constant_0 #(.DATA_WIDTH(1)) constant2(
    .ctrl_valid (fork0_outs_0_valid),
    .ctrl_ready (fork0_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant2_outs),
    .outs_valid (constant2_outs_valid),
    .outs_ready (constant2_outs_ready)
  );

  handshake_cmpi_0 #(.DATA_TYPE(8)) cmpi0(
    .lhs (fork1_outs_0),
    .lhs_valid (fork1_outs_0_valid),
    .lhs_ready (fork1_outs_0_ready),
    .rhs (extsi15_outs),
    .rhs_valid (extsi15_outs_valid),
    .rhs_ready (extsi15_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi0_result),
    .result_valid (cmpi0_result_valid),
    .result_ready (cmpi0_result_ready)
  );

  handshake_cmpi_1 #(.DATA_TYPE(8)) cmpi1(
    .lhs (fork1_outs_1),
    .lhs_valid (fork1_outs_1_valid),
    .lhs_ready (fork1_outs_1_ready),
    .rhs (extsi16_outs),
    .rhs_valid (extsi16_outs_valid),
    .rhs_ready (extsi16_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi1_result),
    .result_valid (cmpi1_result_valid),
    .result_ready (cmpi1_result_ready)
  );

  fork_type #(.SIZE(5), .DATA_TYPE(1)) fork3(
    .ins (cmpi1_result),
    .ins_valid (cmpi1_result_valid),
    .ins_ready (cmpi1_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork3_outs_4, fork3_outs_3, fork3_outs_2, fork3_outs_1, fork3_outs_0}),
    .outs_valid ({fork3_outs_4_valid, fork3_outs_3_valid, fork3_outs_2_valid, fork3_outs_1_valid, fork3_outs_0_valid}),
    .outs_ready ({fork3_outs_4_ready, fork3_outs_3_ready, fork3_outs_2_ready, fork3_outs_1_ready, fork3_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(8)) cond_br3(
    .condition (fork3_outs_0),
    .condition_valid (fork3_outs_0_valid),
    .condition_ready (fork3_outs_0_ready),
    .data (dividend),
    .data_valid (dividend_valid),
    .data_ready (dividend_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br3_trueOut),
    .trueOut_valid (cond_br3_trueOut_valid),
    .trueOut_ready (cond_br3_trueOut_ready),
    .falseOut (cond_br3_falseOut),
    .falseOut_valid (cond_br3_falseOut_valid),
    .falseOut_ready (cond_br3_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink0(
    .ins (cond_br3_falseOut),
    .ins_valid (cond_br3_falseOut_valid),
    .ins_ready (cond_br3_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(8)) cond_br4(
    .condition (fork3_outs_4),
    .condition_valid (fork3_outs_4_valid),
    .condition_ready (fork3_outs_4_ready),
    .data (fork1_outs_2),
    .data_valid (fork1_outs_2_valid),
    .data_ready (fork1_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br4_trueOut),
    .trueOut_valid (cond_br4_trueOut_valid),
    .trueOut_ready (cond_br4_trueOut_ready),
    .falseOut (cond_br4_falseOut),
    .falseOut_valid (cond_br4_falseOut_valid),
    .falseOut_ready (cond_br4_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink1(
    .ins (cond_br4_falseOut),
    .ins_valid (cond_br4_falseOut_valid),
    .ins_ready (cond_br4_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br_dataless cond_br5(
    .condition (fork3_outs_1),
    .condition_valid (fork3_outs_1_valid),
    .condition_ready (fork3_outs_1_ready),
    .data_valid (fork0_outs_2_valid),
    .data_ready (fork0_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br5_trueOut_valid),
    .trueOut_ready (cond_br5_trueOut_ready),
    .falseOut_valid (cond_br5_falseOut_valid),
    .falseOut_ready (cond_br5_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(1)) cond_br6(
    .condition (fork3_outs_3),
    .condition_valid (fork3_outs_3_valid),
    .condition_ready (fork3_outs_3_ready),
    .data (constant2_outs),
    .data_valid (constant2_outs_valid),
    .data_ready (constant2_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br6_trueOut),
    .trueOut_valid (cond_br6_trueOut_valid),
    .trueOut_ready (cond_br6_trueOut_ready),
    .falseOut (cond_br6_falseOut),
    .falseOut_valid (cond_br6_falseOut_valid),
    .falseOut_ready (cond_br6_falseOut_ready)
  );

  sink #(.DATA_TYPE(1)) sink2(
    .ins (cond_br6_trueOut),
    .ins_valid (cond_br6_trueOut_valid),
    .ins_ready (cond_br6_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(1)) cond_br7(
    .condition (fork3_outs_2),
    .condition_valid (fork3_outs_2_valid),
    .condition_ready (fork3_outs_2_ready),
    .data (cmpi0_result),
    .data_valid (cmpi0_result_valid),
    .data_ready (cmpi0_result_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br7_trueOut),
    .trueOut_valid (cond_br7_trueOut_valid),
    .trueOut_ready (cond_br7_trueOut_ready),
    .falseOut (cond_br7_falseOut),
    .falseOut_valid (cond_br7_falseOut_valid),
    .falseOut_ready (cond_br7_falseOut_ready)
  );

  sink #(.DATA_TYPE(1)) sink3(
    .ins (cond_br7_trueOut),
    .ins_valid (cond_br7_trueOut_valid),
    .ins_ready (cond_br7_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(8)) buffer0(
    .ins (cond_br3_trueOut),
    .ins_valid (cond_br3_trueOut_valid),
    .ins_ready (cond_br3_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer0_outs),
    .outs_valid (buffer0_outs_valid),
    .outs_ready (buffer0_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer1(
    .ins (buffer0_outs),
    .ins_valid (buffer0_outs_valid),
    .ins_ready (buffer0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer1_outs),
    .outs_valid (buffer1_outs_valid),
    .outs_ready (buffer1_outs_ready)
  );

  fork_type #(.SIZE(4), .DATA_TYPE(8)) fork4(
    .ins (buffer1_outs),
    .ins_valid (buffer1_outs_valid),
    .ins_ready (buffer1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork4_outs_3, fork4_outs_2, fork4_outs_1, fork4_outs_0}),
    .outs_valid ({fork4_outs_3_valid, fork4_outs_2_valid, fork4_outs_1_valid, fork4_outs_0_valid}),
    .outs_ready ({fork4_outs_3_ready, fork4_outs_2_ready, fork4_outs_1_ready, fork4_outs_0_ready})
  );

  oehb #(.DATA_TYPE(8)) buffer2(
    .ins (cond_br4_trueOut),
    .ins_valid (cond_br4_trueOut_valid),
    .ins_ready (cond_br4_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer2_outs),
    .outs_valid (buffer2_outs_valid),
    .outs_ready (buffer2_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer3(
    .ins (buffer2_outs),
    .ins_valid (buffer2_outs_valid),
    .ins_ready (buffer2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer3_outs),
    .outs_valid (buffer3_outs_valid),
    .outs_ready (buffer3_outs_ready)
  );

  fork_type #(.SIZE(4), .DATA_TYPE(8)) fork5(
    .ins (buffer3_outs),
    .ins_valid (buffer3_outs_valid),
    .ins_ready (buffer3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork5_outs_3, fork5_outs_2, fork5_outs_1, fork5_outs_0}),
    .outs_valid ({fork5_outs_3_valid, fork5_outs_2_valid, fork5_outs_1_valid, fork5_outs_0_valid}),
    .outs_ready ({fork5_outs_3_ready, fork5_outs_2_ready, fork5_outs_1_ready, fork5_outs_0_ready})
  );

  oehb_dataless buffer4(
    .ins_valid (cond_br5_trueOut_valid),
    .ins_ready (cond_br5_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer4_outs_valid),
    .outs_ready (buffer4_outs_ready)
  );

  tehb_dataless buffer5(
    .ins_valid (buffer4_outs_valid),
    .ins_ready (buffer4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer5_outs_valid),
    .outs_ready (buffer5_outs_ready)
  );

  fork_dataless #(.SIZE(2)) fork6(
    .ins_valid (buffer5_outs_valid),
    .ins_ready (buffer5_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork6_outs_1_valid, fork6_outs_0_valid}),
    .outs_ready ({fork6_outs_1_ready, fork6_outs_0_ready})
  );

  source source1(
    .clk (clk),
    .rst (rst),
    .outs_valid (source1_outs_valid),
    .outs_ready (source1_outs_ready)
  );

  handshake_constant_1 #(.DATA_WIDTH(2)) constant3(
    .ctrl_valid (source1_outs_valid),
    .ctrl_ready (source1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant3_outs),
    .outs_valid (constant3_outs_valid),
    .outs_ready (constant3_outs_ready)
  );

  extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(8)) extsi17(
    .ins (constant3_outs),
    .ins_valid (constant3_outs_valid),
    .ins_ready (constant3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi17_outs),
    .outs_valid (extsi17_outs_valid),
    .outs_ready (extsi17_outs_ready)
  );

  source source2(
    .clk (clk),
    .rst (rst),
    .outs_valid (source2_outs_valid),
    .outs_ready (source2_outs_ready)
  );

  handshake_constant_2 #(.DATA_WIDTH(32)) constant7(
    .ctrl_valid (source2_outs_valid),
    .ctrl_ready (source2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant7_outs),
    .outs_valid (constant7_outs_valid),
    .outs_ready (constant7_outs_ready)
  );

  trunci #(.INPUT_TYPE(32), .OUTPUT_TYPE(8)) trunci5(
    .ins (constant7_outs),
    .ins_valid (constant7_outs_valid),
    .ins_ready (constant7_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci5_outs),
    .outs_valid (trunci5_outs_valid),
    .outs_ready (trunci5_outs_ready)
  );

  handshake_constant_0 #(.DATA_WIDTH(1)) constant4(
    .ctrl_valid (fork6_outs_0_valid),
    .ctrl_ready (fork6_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant4_outs),
    .outs_valid (constant4_outs_valid),
    .outs_ready (constant4_outs_ready)
  );

  source source3(
    .clk (clk),
    .rst (rst),
    .outs_valid (source3_outs_valid),
    .outs_ready (source3_outs_ready)
  );

  handshake_constant_0 #(.DATA_WIDTH(1)) constant5(
    .ctrl_valid (source3_outs_valid),
    .ctrl_ready (source3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant5_outs),
    .outs_valid (constant5_outs_valid),
    .outs_ready (constant5_outs_ready)
  );

  fork_type #(.SIZE(6), .DATA_TYPE(1)) fork7(
    .ins (constant5_outs),
    .ins_valid (constant5_outs_valid),
    .ins_ready (constant5_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork7_outs_5, fork7_outs_4, fork7_outs_3, fork7_outs_2, fork7_outs_1, fork7_outs_0}),
    .outs_valid ({fork7_outs_5_valid, fork7_outs_4_valid, fork7_outs_3_valid, fork7_outs_2_valid, fork7_outs_1_valid, fork7_outs_0_valid}),
    .outs_ready ({fork7_outs_5_ready, fork7_outs_4_ready, fork7_outs_3_ready, fork7_outs_2_ready, fork7_outs_1_ready, fork7_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi18(
    .ins (fork7_outs_0),
    .ins_valid (fork7_outs_0_valid),
    .ins_ready (fork7_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi18_outs),
    .outs_valid (extsi18_outs_valid),
    .outs_ready (extsi18_outs_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi19(
    .ins (fork7_outs_1),
    .ins_valid (fork7_outs_1_valid),
    .ins_ready (fork7_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi19_outs),
    .outs_valid (extsi19_outs_valid),
    .outs_ready (extsi19_outs_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi20(
    .ins (fork7_outs_2),
    .ins_valid (fork7_outs_2_valid),
    .ins_ready (fork7_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi20_outs),
    .outs_valid (extsi20_outs_valid),
    .outs_ready (extsi20_outs_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi21(
    .ins (fork7_outs_3),
    .ins_valid (fork7_outs_3_valid),
    .ins_ready (fork7_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi21_outs),
    .outs_valid (extsi21_outs_valid),
    .outs_ready (extsi21_outs_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi22(
    .ins (fork7_outs_4),
    .ins_valid (fork7_outs_4_valid),
    .ins_ready (fork7_outs_4_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi22_outs),
    .outs_valid (extsi22_outs_valid),
    .outs_ready (extsi22_outs_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi23(
    .ins (fork7_outs_5),
    .ins_valid (fork7_outs_5_valid),
    .ins_ready (fork7_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi23_outs),
    .outs_valid (extsi23_outs_valid),
    .outs_ready (extsi23_outs_ready)
  );

  handshake_cmpi_2 #(.DATA_TYPE(8)) cmpi2(
    .lhs (fork4_outs_2),
    .lhs_valid (fork4_outs_2_valid),
    .lhs_ready (fork4_outs_2_ready),
    .rhs (extsi22_outs),
    .rhs_valid (extsi22_outs_valid),
    .rhs_ready (extsi22_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi2_result),
    .result_valid (cmpi2_result_valid),
    .result_ready (cmpi2_result_ready)
  );

  handshake_cmpi_2 #(.DATA_TYPE(8)) cmpi3(
    .lhs (fork5_outs_3),
    .lhs_valid (fork5_outs_3_valid),
    .lhs_ready (fork5_outs_3_ready),
    .rhs (extsi21_outs),
    .rhs_valid (extsi21_outs_valid),
    .rhs_ready (extsi21_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi3_result),
    .result_valid (cmpi3_result_valid),
    .result_ready (cmpi3_result_ready)
  );

  xori #(.DATA_TYPE(1)) xori0(
    .lhs (cmpi2_result),
    .lhs_valid (cmpi2_result_valid),
    .lhs_ready (cmpi2_result_ready),
    .rhs (cmpi3_result),
    .rhs_valid (cmpi3_result_valid),
    .rhs_ready (cmpi3_result_ready),
    .clk (clk),
    .rst (rst),
    .result (xori0_result),
    .result_valid (xori0_result_valid),
    .result_ready (xori0_result_ready)
  );

  selector #(.DATA_TYPE(8)) select0(
    .condition (xori0_result),
    .condition_valid (xori0_result_valid),
    .condition_ready (xori0_result_ready),
    .trueValue (trunci5_outs),
    .trueValue_valid (trunci5_outs_valid),
    .trueValue_ready (trunci5_outs_ready),
    .falseValue (extsi17_outs),
    .falseValue_valid (extsi17_outs_valid),
    .falseValue_ready (extsi17_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (select0_result),
    .result_valid (select0_result_valid),
    .result_ready (select0_result_ready)
  );

  handshake_cmpi_3 #(.DATA_TYPE(8)) cmpi4(
    .lhs (fork4_outs_3),
    .lhs_valid (fork4_outs_3_valid),
    .lhs_ready (fork4_outs_3_ready),
    .rhs (extsi23_outs),
    .rhs_valid (extsi23_outs_valid),
    .rhs_ready (extsi23_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi4_result),
    .result_valid (cmpi4_result_valid),
    .result_ready (cmpi4_result_ready)
  );

  subi #(.DATA_TYPE(8)) subi4(
    .lhs (extsi18_outs),
    .lhs_valid (extsi18_outs_valid),
    .lhs_ready (extsi18_outs_ready),
    .rhs (fork4_outs_0),
    .rhs_valid (fork4_outs_0_valid),
    .rhs_ready (fork4_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .result (subi4_result),
    .result_valid (subi4_result_valid),
    .result_ready (subi4_result_ready)
  );

  selector #(.DATA_TYPE(8)) select2(
    .condition (cmpi4_result),
    .condition_valid (cmpi4_result_valid),
    .condition_ready (cmpi4_result_ready),
    .trueValue (fork4_outs_1),
    .trueValue_valid (fork4_outs_1_valid),
    .trueValue_ready (fork4_outs_1_ready),
    .falseValue (subi4_result),
    .falseValue_valid (subi4_result_valid),
    .falseValue_ready (subi4_result_ready),
    .clk (clk),
    .rst (rst),
    .result (select2_result),
    .result_valid (select2_result_valid),
    .result_ready (select2_result_ready)
  );

  handshake_cmpi_3 #(.DATA_TYPE(8)) cmpi5(
    .lhs (fork5_outs_2),
    .lhs_valid (fork5_outs_2_valid),
    .lhs_ready (fork5_outs_2_ready),
    .rhs (extsi20_outs),
    .rhs_valid (extsi20_outs_valid),
    .rhs_ready (extsi20_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi5_result),
    .result_valid (cmpi5_result_valid),
    .result_ready (cmpi5_result_ready)
  );

  subi #(.DATA_TYPE(8)) subi5(
    .lhs (extsi19_outs),
    .lhs_valid (extsi19_outs_valid),
    .lhs_ready (extsi19_outs_ready),
    .rhs (fork5_outs_0),
    .rhs_valid (fork5_outs_0_valid),
    .rhs_ready (fork5_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .result (subi5_result),
    .result_valid (subi5_result_valid),
    .result_ready (subi5_result_ready)
  );

  selector #(.DATA_TYPE(8)) select3(
    .condition (cmpi5_result),
    .condition_valid (cmpi5_result_valid),
    .condition_ready (cmpi5_result_ready),
    .trueValue (fork5_outs_1),
    .trueValue_valid (fork5_outs_1_valid),
    .trueValue_ready (fork5_outs_1_ready),
    .falseValue (subi5_result),
    .falseValue_valid (subi5_result_valid),
    .falseValue_ready (subi5_result_ready),
    .clk (clk),
    .rst (rst),
    .result (select3_result),
    .result_valid (select3_result_valid),
    .result_ready (select3_result_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi24(
    .ins (constant4_outs),
    .ins_valid (constant4_outs_valid),
    .ins_ready (constant4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi24_outs),
    .outs_valid (extsi24_outs_valid),
    .outs_ready (extsi24_outs_ready)
  );

  mux #(.SIZE(2), .DATA_TYPE(8), .SELECT_TYPE(1)) mux0(
    .index (fork10_outs_1),
    .index_valid (fork10_outs_1_valid),
    .index_ready (fork10_outs_1_ready),
    .ins ({addi0_result, extsi24_outs}),
    .ins_valid ({addi0_result_valid, extsi24_outs_valid}),
    .ins_ready ({addi0_result_ready, extsi24_outs_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux0_outs),
    .outs_valid (mux0_outs_valid),
    .outs_ready (mux0_outs_ready)
  );

  mux #(.SIZE(2), .DATA_TYPE(8), .SELECT_TYPE(1)) mux1(
    .index (fork10_outs_2),
    .index_valid (fork10_outs_2_valid),
    .index_ready (fork10_outs_2_ready),
    .ins ({subi2_result, select2_result}),
    .ins_valid ({subi2_result_valid, select2_result_valid}),
    .ins_ready ({subi2_result_ready, select2_result_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux1_outs),
    .outs_valid (mux1_outs_valid),
    .outs_ready (mux1_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer8(
    .ins (mux1_outs),
    .ins_valid (mux1_outs_valid),
    .ins_ready (mux1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer8_outs),
    .outs_valid (buffer8_outs_valid),
    .outs_ready (buffer8_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer9(
    .ins (buffer8_outs),
    .ins_valid (buffer8_outs_valid),
    .ins_ready (buffer8_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer9_outs),
    .outs_valid (buffer9_outs_valid),
    .outs_ready (buffer9_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(8)) fork8(
    .ins (buffer9_outs),
    .ins_valid (buffer9_outs_valid),
    .ins_ready (buffer9_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork8_outs_1, fork8_outs_0}),
    .outs_valid ({fork8_outs_1_valid, fork8_outs_0_valid}),
    .outs_ready ({fork8_outs_1_ready, fork8_outs_0_ready})
  );

  mux #(.SIZE(2), .DATA_TYPE(8), .SELECT_TYPE(1)) mux2(
    .index (fork10_outs_3),
    .index_valid (fork10_outs_3_valid),
    .index_ready (fork10_outs_3_ready),
    .ins ({buffer21_outs, select0_result}),
    .ins_valid ({buffer21_outs_valid, select0_result_valid}),
    .ins_ready ({buffer21_outs_ready, select0_result_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux2_outs),
    .outs_valid (mux2_outs_valid),
    .outs_ready (mux2_outs_ready)
  );

  mux #(.SIZE(2), .DATA_TYPE(8), .SELECT_TYPE(1)) mux3(
    .index (fork10_outs_0),
    .index_valid (fork10_outs_0_valid),
    .index_ready (fork10_outs_0_ready),
    .ins ({fork12_outs_1, select3_result}),
    .ins_valid ({fork12_outs_1_valid, select3_result_valid}),
    .ins_ready ({fork12_outs_1_ready, select3_result_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux3_outs),
    .outs_valid (mux3_outs_valid),
    .outs_ready (mux3_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer12(
    .ins (mux3_outs),
    .ins_valid (mux3_outs_valid),
    .ins_ready (mux3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer12_outs),
    .outs_valid (buffer12_outs_valid),
    .outs_ready (buffer12_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer13(
    .ins (buffer12_outs),
    .ins_valid (buffer12_outs_valid),
    .ins_ready (buffer12_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer13_outs),
    .outs_valid (buffer13_outs_valid),
    .outs_ready (buffer13_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(8)) fork9(
    .ins (buffer13_outs),
    .ins_valid (buffer13_outs_valid),
    .ins_ready (buffer13_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork9_outs_1, fork9_outs_0}),
    .outs_valid ({fork9_outs_1_valid, fork9_outs_0_valid}),
    .outs_ready ({fork9_outs_1_ready, fork9_outs_0_ready})
  );

  control_merge_dataless #(.SIZE(2), .INDEX_TYPE(1)) control_merge1(
    .ins_valid ({buffer25_outs_valid, fork6_outs_1_valid}),
    .ins_ready ({buffer25_outs_ready, fork6_outs_1_ready}),
    .clk (clk),
    .rst (rst),
    .outs_valid (control_merge1_outs_valid),
    .outs_ready (control_merge1_outs_ready),
    .index (control_merge1_index),
    .index_valid (control_merge1_index_valid),
    .index_ready (control_merge1_index_ready)
  );

  fork_type #(.SIZE(4), .DATA_TYPE(1)) fork10(
    .ins (control_merge1_index),
    .ins_valid (control_merge1_index_valid),
    .ins_ready (control_merge1_index_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork10_outs_3, fork10_outs_2, fork10_outs_1, fork10_outs_0}),
    .outs_valid ({fork10_outs_3_valid, fork10_outs_2_valid, fork10_outs_1_valid, fork10_outs_0_valid}),
    .outs_ready ({fork10_outs_3_ready, fork10_outs_2_ready, fork10_outs_1_ready, fork10_outs_0_ready})
  );

  handshake_cmpi_3 #(.DATA_TYPE(8)) cmpi6(
    .lhs (fork8_outs_0),
    .lhs_valid (fork8_outs_0_valid),
    .lhs_ready (fork8_outs_0_ready),
    .rhs (fork9_outs_1),
    .rhs_valid (fork9_outs_1_valid),
    .rhs_ready (fork9_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi6_result),
    .result_valid (cmpi6_result_valid),
    .result_ready (cmpi6_result_ready)
  );

  fork_type #(.SIZE(5), .DATA_TYPE(1)) fork11(
    .ins (cmpi6_result),
    .ins_valid (cmpi6_result_valid),
    .ins_ready (cmpi6_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork11_outs_4, fork11_outs_3, fork11_outs_2, fork11_outs_1, fork11_outs_0}),
    .outs_valid ({fork11_outs_4_valid, fork11_outs_3_valid, fork11_outs_2_valid, fork11_outs_1_valid, fork11_outs_0_valid}),
    .outs_ready ({fork11_outs_4_ready, fork11_outs_3_ready, fork11_outs_2_ready, fork11_outs_1_ready, fork11_outs_0_ready})
  );

  oehb #(.DATA_TYPE(8)) buffer6(
    .ins (mux0_outs),
    .ins_valid (mux0_outs_valid),
    .ins_ready (mux0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer6_outs),
    .outs_valid (buffer6_outs_valid),
    .outs_ready (buffer6_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer7(
    .ins (buffer6_outs),
    .ins_valid (buffer6_outs_valid),
    .ins_ready (buffer6_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer7_outs),
    .outs_valid (buffer7_outs_valid),
    .outs_ready (buffer7_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br8(
    .condition (fork11_outs_1),
    .condition_valid (fork11_outs_1_valid),
    .condition_ready (fork11_outs_1_ready),
    .data (buffer7_outs),
    .data_valid (buffer7_outs_valid),
    .data_ready (buffer7_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br8_trueOut),
    .trueOut_valid (cond_br8_trueOut_valid),
    .trueOut_ready (cond_br8_trueOut_ready),
    .falseOut (cond_br8_falseOut),
    .falseOut_valid (cond_br8_falseOut_valid),
    .falseOut_ready (cond_br8_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br9(
    .condition (fork11_outs_2),
    .condition_valid (fork11_outs_2_valid),
    .condition_ready (fork11_outs_2_ready),
    .data (fork8_outs_1),
    .data_valid (fork8_outs_1_valid),
    .data_ready (fork8_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br9_trueOut),
    .trueOut_valid (cond_br9_trueOut_valid),
    .trueOut_ready (cond_br9_trueOut_ready),
    .falseOut (cond_br9_falseOut),
    .falseOut_valid (cond_br9_falseOut_valid),
    .falseOut_ready (cond_br9_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink5(
    .ins (cond_br9_falseOut),
    .ins_valid (cond_br9_falseOut_valid),
    .ins_ready (cond_br9_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(8)) buffer10(
    .ins (mux2_outs),
    .ins_valid (mux2_outs_valid),
    .ins_ready (mux2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer10_outs),
    .outs_valid (buffer10_outs_valid),
    .outs_ready (buffer10_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer11(
    .ins (buffer10_outs),
    .ins_valid (buffer10_outs_valid),
    .ins_ready (buffer10_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer11_outs),
    .outs_valid (buffer11_outs_valid),
    .outs_ready (buffer11_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br10(
    .condition (fork11_outs_3),
    .condition_valid (fork11_outs_3_valid),
    .condition_ready (fork11_outs_3_ready),
    .data (buffer11_outs),
    .data_valid (buffer11_outs_valid),
    .data_ready (buffer11_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br10_trueOut),
    .trueOut_valid (cond_br10_trueOut_valid),
    .trueOut_ready (cond_br10_trueOut_ready),
    .falseOut (cond_br10_falseOut),
    .falseOut_valid (cond_br10_falseOut_valid),
    .falseOut_ready (cond_br10_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br11(
    .condition (fork11_outs_0),
    .condition_valid (fork11_outs_0_valid),
    .condition_ready (fork11_outs_0_ready),
    .data (fork9_outs_0),
    .data_valid (fork9_outs_0_valid),
    .data_ready (fork9_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br11_trueOut),
    .trueOut_valid (cond_br11_trueOut_valid),
    .trueOut_ready (cond_br11_trueOut_ready),
    .falseOut (cond_br11_falseOut),
    .falseOut_valid (cond_br11_falseOut_valid),
    .falseOut_ready (cond_br11_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink6(
    .ins (cond_br11_falseOut),
    .ins_valid (cond_br11_falseOut_valid),
    .ins_ready (cond_br11_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb_dataless buffer14(
    .ins_valid (control_merge1_outs_valid),
    .ins_ready (control_merge1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer14_outs_valid),
    .outs_ready (buffer14_outs_ready)
  );

  tehb_dataless buffer15(
    .ins_valid (buffer14_outs_valid),
    .ins_ready (buffer14_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer15_outs_valid),
    .outs_ready (buffer15_outs_ready)
  );

  cond_br_dataless cond_br12(
    .condition (fork11_outs_4),
    .condition_valid (fork11_outs_4_valid),
    .condition_ready (fork11_outs_4_ready),
    .data_valid (buffer15_outs_valid),
    .data_ready (buffer15_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br12_trueOut_valid),
    .trueOut_ready (cond_br12_trueOut_ready),
    .falseOut_valid (cond_br12_falseOut_valid),
    .falseOut_ready (cond_br12_falseOut_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer22(
    .ins (cond_br11_trueOut),
    .ins_valid (cond_br11_trueOut_valid),
    .ins_ready (cond_br11_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer22_outs),
    .outs_valid (buffer22_outs_valid),
    .outs_ready (buffer22_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer23(
    .ins (buffer22_outs),
    .ins_valid (buffer22_outs_valid),
    .ins_ready (buffer22_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer23_outs),
    .outs_valid (buffer23_outs_valid),
    .outs_ready (buffer23_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(8)) fork12(
    .ins (buffer23_outs),
    .ins_valid (buffer23_outs_valid),
    .ins_ready (buffer23_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork12_outs_1, fork12_outs_0}),
    .outs_valid ({fork12_outs_1_valid, fork12_outs_0_valid}),
    .outs_ready ({fork12_outs_1_ready, fork12_outs_0_ready})
  );

  source source4(
    .clk (clk),
    .rst (rst),
    .outs_valid (source4_outs_valid),
    .outs_ready (source4_outs_ready)
  );

  handshake_constant_1 #(.DATA_WIDTH(2)) constant14(
    .ctrl_valid (source4_outs_valid),
    .ctrl_ready (source4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant14_outs),
    .outs_valid (constant14_outs_valid),
    .outs_ready (constant14_outs_ready)
  );

  extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(8)) extsi13(
    .ins (constant14_outs),
    .ins_valid (constant14_outs_valid),
    .ins_ready (constant14_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi13_outs),
    .outs_valid (extsi13_outs_valid),
    .outs_ready (extsi13_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer18(
    .ins (cond_br9_trueOut),
    .ins_valid (cond_br9_trueOut_valid),
    .ins_ready (cond_br9_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer18_outs),
    .outs_valid (buffer18_outs_valid),
    .outs_ready (buffer18_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer19(
    .ins (buffer18_outs),
    .ins_valid (buffer18_outs_valid),
    .ins_ready (buffer18_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer19_outs),
    .outs_valid (buffer19_outs_valid),
    .outs_ready (buffer19_outs_ready)
  );

  subi #(.DATA_TYPE(8)) subi2(
    .lhs (buffer19_outs),
    .lhs_valid (buffer19_outs_valid),
    .lhs_ready (buffer19_outs_ready),
    .rhs (fork12_outs_0),
    .rhs_valid (fork12_outs_0_valid),
    .rhs_ready (fork12_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .result (subi2_result),
    .result_valid (subi2_result_valid),
    .result_ready (subi2_result_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer16(
    .ins (cond_br8_trueOut),
    .ins_valid (cond_br8_trueOut_valid),
    .ins_ready (cond_br8_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer16_outs),
    .outs_valid (buffer16_outs_valid),
    .outs_ready (buffer16_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer17(
    .ins (buffer16_outs),
    .ins_valid (buffer16_outs_valid),
    .ins_ready (buffer16_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer17_outs),
    .outs_valid (buffer17_outs_valid),
    .outs_ready (buffer17_outs_ready)
  );

  addi #(.DATA_TYPE(8)) addi0(
    .lhs (buffer17_outs),
    .lhs_valid (buffer17_outs_valid),
    .lhs_ready (buffer17_outs_ready),
    .rhs (extsi13_outs),
    .rhs_valid (extsi13_outs_valid),
    .rhs_ready (extsi13_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi0_result),
    .result_valid (addi0_result_valid),
    .result_ready (addi0_result_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer20(
    .ins (cond_br10_trueOut),
    .ins_valid (cond_br10_trueOut_valid),
    .ins_ready (cond_br10_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer20_outs),
    .outs_valid (buffer20_outs_valid),
    .outs_ready (buffer20_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer21(
    .ins (buffer20_outs),
    .ins_valid (buffer20_outs_valid),
    .ins_ready (buffer20_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer21_outs),
    .outs_valid (buffer21_outs_valid),
    .outs_ready (buffer21_outs_ready)
  );

  oehb_dataless buffer24(
    .ins_valid (cond_br12_trueOut_valid),
    .ins_ready (cond_br12_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer24_outs_valid),
    .outs_ready (buffer24_outs_ready)
  );

  tehb_dataless buffer25(
    .ins_valid (buffer24_outs_valid),
    .ins_ready (buffer24_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer25_outs_valid),
    .outs_ready (buffer25_outs_ready)
  );

  source source5(
    .clk (clk),
    .rst (rst),
    .outs_valid (source5_outs_valid),
    .outs_ready (source5_outs_ready)
  );

  handshake_constant_2 #(.DATA_WIDTH(32)) constant11(
    .ctrl_valid (source5_outs_valid),
    .ctrl_ready (source5_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant11_outs),
    .outs_valid (constant11_outs_valid),
    .outs_ready (constant11_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer26(
    .ins (cond_br10_falseOut),
    .ins_valid (cond_br10_falseOut_valid),
    .ins_ready (cond_br10_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer26_outs),
    .outs_valid (buffer26_outs_valid),
    .outs_ready (buffer26_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer27(
    .ins (buffer26_outs),
    .ins_valid (buffer26_outs_valid),
    .ins_ready (buffer26_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer27_outs),
    .outs_valid (buffer27_outs_valid),
    .outs_ready (buffer27_outs_ready)
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(32)) extsi5(
    .ins (buffer27_outs),
    .ins_valid (buffer27_outs_valid),
    .ins_ready (buffer27_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi5_outs),
    .outs_valid (extsi5_outs_valid),
    .outs_ready (extsi5_outs_ready)
  );

  handshake_cmpi_4 #(.DATA_TYPE(32)) cmpi7(
    .lhs (extsi5_outs),
    .lhs_valid (extsi5_outs_valid),
    .lhs_ready (extsi5_outs_ready),
    .rhs (constant11_outs),
    .rhs_valid (constant11_outs_valid),
    .rhs_ready (constant11_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi7_result),
    .result_valid (cmpi7_result_valid),
    .result_ready (cmpi7_result_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(1)) fork13(
    .ins (cmpi7_result),
    .ins_valid (cmpi7_result_valid),
    .ins_ready (cmpi7_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork13_outs_1, fork13_outs_0}),
    .outs_valid ({fork13_outs_1_valid, fork13_outs_0_valid}),
    .outs_ready ({fork13_outs_1_ready, fork13_outs_0_ready})
  );

  oehb #(.DATA_TYPE(8)) buffer28(
    .ins (cond_br8_falseOut),
    .ins_valid (cond_br8_falseOut_valid),
    .ins_ready (cond_br8_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer28_outs),
    .outs_valid (buffer28_outs_valid),
    .outs_ready (buffer28_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer29(
    .ins (buffer28_outs),
    .ins_valid (buffer28_outs_valid),
    .ins_ready (buffer28_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer29_outs),
    .outs_valid (buffer29_outs_valid),
    .outs_ready (buffer29_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br13(
    .condition (fork13_outs_1),
    .condition_valid (fork13_outs_1_valid),
    .condition_ready (fork13_outs_1_ready),
    .data (buffer29_outs),
    .data_valid (buffer29_outs_valid),
    .data_ready (buffer29_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br13_trueOut),
    .trueOut_valid (cond_br13_trueOut_valid),
    .trueOut_ready (cond_br13_trueOut_ready),
    .falseOut (cond_br13_falseOut),
    .falseOut_valid (cond_br13_falseOut_valid),
    .falseOut_ready (cond_br13_falseOut_ready)
  );

  oehb_dataless buffer30(
    .ins_valid (cond_br12_falseOut_valid),
    .ins_ready (cond_br12_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer30_outs_valid),
    .outs_ready (buffer30_outs_ready)
  );

  tehb_dataless buffer31(
    .ins_valid (buffer30_outs_valid),
    .ins_ready (buffer30_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer31_outs_valid),
    .outs_ready (buffer31_outs_ready)
  );

  cond_br_dataless cond_br14(
    .condition (fork13_outs_0),
    .condition_valid (fork13_outs_0_valid),
    .condition_ready (fork13_outs_0_ready),
    .data_valid (buffer31_outs_valid),
    .data_ready (buffer31_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br14_trueOut_valid),
    .trueOut_ready (cond_br14_trueOut_ready),
    .falseOut_valid (cond_br14_falseOut_valid),
    .falseOut_ready (cond_br14_falseOut_ready)
  );

  source source6(
    .clk (clk),
    .rst (rst),
    .outs_valid (source6_outs_valid),
    .outs_ready (source6_outs_ready)
  );

  handshake_constant_0 #(.DATA_WIDTH(1)) constant15(
    .ctrl_valid (source6_outs_valid),
    .ctrl_ready (source6_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant15_outs),
    .outs_valid (constant15_outs_valid),
    .outs_ready (constant15_outs_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi25(
    .ins (constant15_outs),
    .ins_valid (constant15_outs_valid),
    .ins_ready (constant15_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi25_outs),
    .outs_valid (extsi25_outs_valid),
    .outs_ready (extsi25_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer32(
    .ins (cond_br13_trueOut),
    .ins_valid (cond_br13_trueOut_valid),
    .ins_ready (cond_br13_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer32_outs),
    .outs_valid (buffer32_outs_valid),
    .outs_ready (buffer32_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer33(
    .ins (buffer32_outs),
    .ins_valid (buffer32_outs_valid),
    .ins_ready (buffer32_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer33_outs),
    .outs_valid (buffer33_outs_valid),
    .outs_ready (buffer33_outs_ready)
  );

  subi #(.DATA_TYPE(8)) subi3(
    .lhs (extsi25_outs),
    .lhs_valid (extsi25_outs_valid),
    .lhs_ready (extsi25_outs_ready),
    .rhs (buffer33_outs),
    .rhs_valid (buffer33_outs_valid),
    .rhs_ready (buffer33_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (subi3_result),
    .result_valid (subi3_result_valid),
    .result_ready (subi3_result_ready)
  );

  oehb_dataless buffer34(
    .ins_valid (cond_br14_trueOut_valid),
    .ins_ready (cond_br14_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer34_outs_valid),
    .outs_ready (buffer34_outs_ready)
  );

  tehb_dataless buffer35(
    .ins_valid (buffer34_outs_valid),
    .ins_ready (buffer34_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer35_outs_valid),
    .outs_ready (buffer35_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer36(
    .ins (cond_br13_falseOut),
    .ins_valid (cond_br13_falseOut_valid),
    .ins_ready (cond_br13_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer36_outs),
    .outs_valid (buffer36_outs_valid),
    .outs_ready (buffer36_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer37(
    .ins (buffer36_outs),
    .ins_valid (buffer36_outs_valid),
    .ins_ready (buffer36_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer37_outs),
    .outs_valid (buffer37_outs_valid),
    .outs_ready (buffer37_outs_ready)
  );

  oehb_dataless buffer38(
    .ins_valid (cond_br14_falseOut_valid),
    .ins_ready (cond_br14_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer38_outs_valid),
    .outs_ready (buffer38_outs_ready)
  );

  tehb_dataless buffer39(
    .ins_valid (buffer38_outs_valid),
    .ins_ready (buffer38_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer39_outs_valid),
    .outs_ready (buffer39_outs_ready)
  );

  mux #(.SIZE(2), .DATA_TYPE(8), .SELECT_TYPE(1)) mux4(
    .index (control_merge6_index),
    .index_valid (control_merge6_index_valid),
    .index_ready (control_merge6_index_ready),
    .ins ({buffer37_outs, subi3_result}),
    .ins_valid ({buffer37_outs_valid, subi3_result_valid}),
    .ins_ready ({buffer37_outs_ready, subi3_result_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux4_outs),
    .outs_valid (mux4_outs_valid),
    .outs_ready (mux4_outs_ready)
  );

  control_merge_dataless #(.SIZE(2), .INDEX_TYPE(1)) control_merge6(
    .ins_valid ({buffer39_outs_valid, buffer35_outs_valid}),
    .ins_ready ({buffer39_outs_ready, buffer35_outs_ready}),
    .clk (clk),
    .rst (rst),
    .outs_valid (control_merge6_outs_valid),
    .outs_ready (control_merge6_outs_ready),
    .index (control_merge6_index),
    .index_valid (control_merge6_index_valid),
    .index_ready (control_merge6_index_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer40(
    .ins (mux4_outs),
    .ins_valid (mux4_outs_valid),
    .ins_ready (mux4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer40_outs),
    .outs_valid (buffer40_outs_valid),
    .outs_ready (buffer40_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer41(
    .ins (buffer40_outs),
    .ins_valid (buffer40_outs_valid),
    .ins_ready (buffer40_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer41_outs),
    .outs_valid (buffer41_outs_valid),
    .outs_ready (buffer41_outs_ready)
  );

  oehb_dataless buffer42(
    .ins_valid (control_merge6_outs_valid),
    .ins_ready (control_merge6_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer42_outs_valid),
    .outs_ready (buffer42_outs_ready)
  );

  tehb_dataless buffer43(
    .ins_valid (buffer42_outs_valid),
    .ins_ready (buffer42_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer43_outs_valid),
    .outs_ready (buffer43_outs_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer44(
    .ins (cond_br6_falseOut),
    .ins_valid (cond_br6_falseOut_valid),
    .ins_ready (cond_br6_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer44_outs),
    .outs_valid (buffer44_outs_valid),
    .outs_ready (buffer44_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer45(
    .ins (buffer44_outs),
    .ins_valid (buffer44_outs_valid),
    .ins_ready (buffer44_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer45_outs),
    .outs_valid (buffer45_outs_valid),
    .outs_ready (buffer45_outs_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi26(
    .ins (buffer45_outs),
    .ins_valid (buffer45_outs_valid),
    .ins_ready (buffer45_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi26_outs),
    .outs_valid (extsi26_outs_valid),
    .outs_ready (extsi26_outs_ready)
  );

  source source7(
    .clk (clk),
    .rst (rst),
    .outs_valid (source7_outs_valid),
    .outs_ready (source7_outs_ready)
  );

  handshake_constant_3 #(.DATA_WIDTH(8)) constant13(
    .ctrl_valid (source7_outs_valid),
    .ctrl_ready (source7_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant13_outs),
    .outs_valid (constant13_outs_valid),
    .outs_ready (constant13_outs_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer46(
    .ins (cond_br7_falseOut),
    .ins_valid (cond_br7_falseOut_valid),
    .ins_ready (cond_br7_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer46_outs),
    .outs_valid (buffer46_outs_valid),
    .outs_ready (buffer46_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer47(
    .ins (buffer46_outs),
    .ins_valid (buffer46_outs_valid),
    .ins_ready (buffer46_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer47_outs),
    .outs_valid (buffer47_outs_valid),
    .outs_ready (buffer47_outs_ready)
  );

  selector #(.DATA_TYPE(8)) select1(
    .condition (buffer47_outs),
    .condition_valid (buffer47_outs_valid),
    .condition_ready (buffer47_outs_ready),
    .trueValue (constant13_outs),
    .trueValue_valid (constant13_outs_valid),
    .trueValue_ready (constant13_outs_ready),
    .falseValue (extsi26_outs),
    .falseValue_valid (extsi26_outs_valid),
    .falseValue_ready (extsi26_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (select1_result),
    .result_valid (select1_result_valid),
    .result_ready (select1_result_ready)
  );

  oehb_dataless buffer48(
    .ins_valid (cond_br5_falseOut_valid),
    .ins_ready (cond_br5_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer48_outs_valid),
    .outs_ready (buffer48_outs_ready)
  );

  tehb_dataless buffer49(
    .ins_valid (buffer48_outs_valid),
    .ins_ready (buffer48_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer49_outs_valid),
    .outs_ready (buffer49_outs_ready)
  );

  mux #(.SIZE(2), .DATA_TYPE(8), .SELECT_TYPE(1)) mux5(
    .index (control_merge8_index),
    .index_valid (control_merge8_index_valid),
    .index_ready (control_merge8_index_ready),
    .ins ({select1_result, buffer41_outs}),
    .ins_valid ({select1_result_valid, buffer41_outs_valid}),
    .ins_ready ({select1_result_ready, buffer41_outs_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux5_outs),
    .outs_valid (mux5_outs_valid),
    .outs_ready (mux5_outs_ready)
  );

  control_merge_dataless #(.SIZE(2), .INDEX_TYPE(1)) control_merge8(
    .ins_valid ({buffer49_outs_valid, buffer43_outs_valid}),
    .ins_ready ({buffer49_outs_ready, buffer43_outs_ready}),
    .clk (clk),
    .rst (rst),
    .outs_valid (control_merge8_outs_valid),
    .outs_ready (control_merge8_outs_ready),
    .index (control_merge8_index),
    .index_valid (control_merge8_index_valid),
    .index_ready (control_merge8_index_ready)
  );

  oehb_dataless buffer52(
    .ins_valid (control_merge8_outs_valid),
    .ins_ready (control_merge8_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer52_outs_valid),
    .outs_ready (buffer52_outs_ready)
  );

  tehb_dataless buffer53(
    .ins_valid (buffer52_outs_valid),
    .ins_ready (buffer52_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer53_outs_valid),
    .outs_ready (buffer53_outs_ready)
  );

  sink_dataless sink12(
    .ins_valid (buffer53_outs_valid),
    .ins_ready (buffer53_outs_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(8)) buffer50(
    .ins (mux5_outs),
    .ins_valid (mux5_outs_valid),
    .ins_ready (mux5_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer50_outs),
    .outs_valid (buffer50_outs_valid),
    .outs_ready (buffer50_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer51(
    .ins (buffer50_outs),
    .ins_valid (buffer50_outs_valid),
    .ins_ready (buffer50_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer51_outs),
    .outs_valid (buffer51_outs_valid),
    .outs_ready (buffer51_outs_ready)
  );

endmodule
