`timescale 1ns/1ns
module tb;
reg [0:0] arg0_valid; // input signal
reg [0:0] out0_ready; // input signal
reg [0:0] rst; // input signal
reg [9:0] arg0; // input signal
wire [0:0] arg0_ready; // output signal
wire [0:0] out0_valid; // output signal
wire [9:0] out0; // output signal
reg clk = 0;
main dut(
.arg0_valid(arg0_valid),
.clk(clk),
.out0_ready(out0_ready),
.rst(rst),
.arg0(arg0),
.arg0_ready(arg0_ready),
.out0_valid(out0_valid),
.out0(out0)
);
always
	 #2 clk = ~clk;
initial begin
$dumpfile("./trace_round_0.vcd");
$dumpvars(0, tb.dut);
arg0_valid <= 1;
out0_ready <= 0;
rst <= 1;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 3;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 1;
rst <= 0;
arg0 <= 1;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 0;
out0_ready <= 0;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 2;
#4;
arg0_valid <= 1;
out0_ready <= 1;
rst <= 0;
arg0 <= 0;
#4;
arg0_valid <= 1;
out0_ready <= 0;
rst <= 0;
arg0 <= 1;
#4;
$finish;
end
endmodule
