module iterative_sqrt(
  input [7:0] n,
  input  n_valid,
  input  start_valid,
  input  clk,
  input  rst,
  input  out0_ready,
  input  end_ready,
  output  n_ready,
  output  start_ready,
  output [7:0] out0,
  output  out0_valid,
  output  end_valid
);
  wire  fork0_outs_0_valid;
  wire  fork0_outs_0_ready;
  wire  fork0_outs_1_valid;
  wire  fork0_outs_1_ready;
  wire  fork0_outs_2_valid;
  wire  fork0_outs_2_ready;
  wire  fork0_outs_3_valid;
  wire  fork0_outs_3_ready;
  wire [7:0] fork1_outs_0;
  wire  fork1_outs_0_valid;
  wire  fork1_outs_0_ready;
  wire [7:0] fork1_outs_1;
  wire  fork1_outs_1_valid;
  wire  fork1_outs_1_ready;
  wire [0:0] constant1_outs;
  wire  constant1_outs_valid;
  wire  constant1_outs_ready;
  wire [0:0] fork2_outs_0;
  wire  fork2_outs_0_valid;
  wire  fork2_outs_0_ready;
  wire [0:0] fork2_outs_1;
  wire  fork2_outs_1_valid;
  wire  fork2_outs_1_ready;
  wire [0:0] constant3_outs;
  wire  constant3_outs_valid;
  wire  constant3_outs_ready;
  wire [7:0] extsi10_outs;
  wire  extsi10_outs_valid;
  wire  extsi10_outs_ready;
  wire [0:0] fork3_outs_0;
  wire  fork3_outs_0_valid;
  wire  fork3_outs_0_ready;
  wire [0:0] fork3_outs_1;
  wire  fork3_outs_1_valid;
  wire  fork3_outs_1_ready;
  wire [7:0] extsi11_outs;
  wire  extsi11_outs_valid;
  wire  extsi11_outs_ready;
  wire [7:0] mux0_outs;
  wire  mux0_outs_valid;
  wire  mux0_outs_ready;
  wire [7:0] buffer0_outs;
  wire  buffer0_outs_valid;
  wire  buffer0_outs_ready;
  wire [7:0] buffer1_outs;
  wire  buffer1_outs_valid;
  wire  buffer1_outs_ready;
  wire [7:0] fork4_outs_0;
  wire  fork4_outs_0_valid;
  wire  fork4_outs_0_ready;
  wire [7:0] fork4_outs_1;
  wire  fork4_outs_1_valid;
  wire  fork4_outs_1_ready;
  wire [7:0] mux1_outs;
  wire  mux1_outs_valid;
  wire  mux1_outs_ready;
  wire [7:0] buffer2_outs;
  wire  buffer2_outs_valid;
  wire  buffer2_outs_ready;
  wire [7:0] buffer3_outs;
  wire  buffer3_outs_valid;
  wire  buffer3_outs_ready;
  wire [7:0] fork5_outs_0;
  wire  fork5_outs_0_valid;
  wire  fork5_outs_0_ready;
  wire [7:0] fork5_outs_1;
  wire  fork5_outs_1_valid;
  wire  fork5_outs_1_ready;
  wire [0:0] mux2_outs;
  wire  mux2_outs_valid;
  wire  mux2_outs_ready;
  wire [7:0] mux3_outs;
  wire  mux3_outs_valid;
  wire  mux3_outs_ready;
  wire [0:0] mux4_outs;
  wire  mux4_outs_valid;
  wire  mux4_outs_ready;
  wire [7:0] mux5_outs;
  wire  mux5_outs_valid;
  wire  mux5_outs_ready;
  wire  control_merge0_outs_valid;
  wire  control_merge0_outs_ready;
  wire [1:0] control_merge0_index;
  wire  control_merge0_index_valid;
  wire  control_merge0_index_ready;
  wire [1:0] fork6_outs_0;
  wire  fork6_outs_0_valid;
  wire  fork6_outs_0_ready;
  wire [1:0] fork6_outs_1;
  wire  fork6_outs_1_valid;
  wire  fork6_outs_1_ready;
  wire [1:0] fork6_outs_2;
  wire  fork6_outs_2_valid;
  wire  fork6_outs_2_ready;
  wire [1:0] fork6_outs_3;
  wire  fork6_outs_3_valid;
  wire  fork6_outs_3_ready;
  wire [1:0] fork6_outs_4;
  wire  fork6_outs_4_valid;
  wire  fork6_outs_4_ready;
  wire [1:0] fork6_outs_5;
  wire  fork6_outs_5_valid;
  wire  fork6_outs_5_ready;
  wire [0:0] cmpi0_result;
  wire  cmpi0_result_valid;
  wire  cmpi0_result_ready;
  wire [0:0] buffer8_outs;
  wire  buffer8_outs_valid;
  wire  buffer8_outs_ready;
  wire [0:0] buffer9_outs;
  wire  buffer9_outs_valid;
  wire  buffer9_outs_ready;
  wire [0:0] andi0_result;
  wire  andi0_result_valid;
  wire  andi0_result_ready;
  wire [0:0] fork7_outs_0;
  wire  fork7_outs_0_valid;
  wire  fork7_outs_0_ready;
  wire [0:0] fork7_outs_1;
  wire  fork7_outs_1_valid;
  wire  fork7_outs_1_ready;
  wire [0:0] fork7_outs_2;
  wire  fork7_outs_2_valid;
  wire  fork7_outs_2_ready;
  wire [0:0] fork7_outs_3;
  wire  fork7_outs_3_valid;
  wire  fork7_outs_3_ready;
  wire [0:0] fork7_outs_4;
  wire  fork7_outs_4_valid;
  wire  fork7_outs_4_ready;
  wire [0:0] fork7_outs_5;
  wire  fork7_outs_5_valid;
  wire  fork7_outs_5_ready;
  wire [7:0] cond_br3_trueOut;
  wire  cond_br3_trueOut_valid;
  wire  cond_br3_trueOut_ready;
  wire [7:0] cond_br3_falseOut;
  wire  cond_br3_falseOut_valid;
  wire  cond_br3_falseOut_ready;
  wire [0:0] buffer4_outs;
  wire  buffer4_outs_valid;
  wire  buffer4_outs_ready;
  wire [0:0] buffer5_outs;
  wire  buffer5_outs_valid;
  wire  buffer5_outs_ready;
  wire [0:0] cond_br4_trueOut;
  wire  cond_br4_trueOut_valid;
  wire  cond_br4_trueOut_ready;
  wire [0:0] cond_br4_falseOut;
  wire  cond_br4_falseOut_valid;
  wire  cond_br4_falseOut_ready;
  wire [7:0] buffer6_outs;
  wire  buffer6_outs_valid;
  wire  buffer6_outs_ready;
  wire [7:0] buffer7_outs;
  wire  buffer7_outs_valid;
  wire  buffer7_outs_ready;
  wire [7:0] cond_br5_trueOut;
  wire  cond_br5_trueOut_valid;
  wire  cond_br5_trueOut_ready;
  wire [7:0] cond_br5_falseOut;
  wire  cond_br5_falseOut_valid;
  wire  cond_br5_falseOut_ready;
  wire [7:0] cond_br6_trueOut;
  wire  cond_br6_trueOut_valid;
  wire  cond_br6_trueOut_ready;
  wire [7:0] cond_br6_falseOut;
  wire  cond_br6_falseOut_valid;
  wire  cond_br6_falseOut_ready;
  wire [7:0] buffer10_outs;
  wire  buffer10_outs_valid;
  wire  buffer10_outs_ready;
  wire [7:0] buffer11_outs;
  wire  buffer11_outs_valid;
  wire  buffer11_outs_ready;
  wire [7:0] cond_br7_trueOut;
  wire  cond_br7_trueOut_valid;
  wire  cond_br7_trueOut_ready;
  wire [7:0] cond_br7_falseOut;
  wire  cond_br7_falseOut_valid;
  wire  cond_br7_falseOut_ready;
  wire  buffer12_outs_valid;
  wire  buffer12_outs_ready;
  wire  buffer13_outs_valid;
  wire  buffer13_outs_ready;
  wire  cond_br8_trueOut_valid;
  wire  cond_br8_trueOut_ready;
  wire  cond_br8_falseOut_valid;
  wire  cond_br8_falseOut_ready;
  wire [7:0] buffer14_outs;
  wire  buffer14_outs_valid;
  wire  buffer14_outs_ready;
  wire [7:0] buffer15_outs;
  wire  buffer15_outs_valid;
  wire  buffer15_outs_ready;
  wire [7:0] fork8_outs_0;
  wire  fork8_outs_0_valid;
  wire  fork8_outs_0_ready;
  wire [7:0] fork8_outs_1;
  wire  fork8_outs_1_valid;
  wire  fork8_outs_1_ready;
  wire [8:0] extsi12_outs;
  wire  extsi12_outs_valid;
  wire  extsi12_outs_ready;
  wire [7:0] buffer20_outs;
  wire  buffer20_outs_valid;
  wire  buffer20_outs_ready;
  wire [7:0] buffer21_outs;
  wire  buffer21_outs_valid;
  wire  buffer21_outs_ready;
  wire [7:0] fork9_outs_0;
  wire  fork9_outs_0_valid;
  wire  fork9_outs_0_ready;
  wire [7:0] fork9_outs_1;
  wire  fork9_outs_1_valid;
  wire  fork9_outs_1_ready;
  wire [8:0] extsi13_outs;
  wire  extsi13_outs_valid;
  wire  extsi13_outs_ready;
  wire [7:0] buffer22_outs;
  wire  buffer22_outs_valid;
  wire  buffer22_outs_ready;
  wire [7:0] buffer23_outs;
  wire  buffer23_outs_valid;
  wire  buffer23_outs_ready;
  wire [7:0] fork10_outs_0;
  wire  fork10_outs_0_valid;
  wire  fork10_outs_0_ready;
  wire [7:0] fork10_outs_1;
  wire  fork10_outs_1_valid;
  wire  fork10_outs_1_ready;
  wire [7:0] fork10_outs_2;
  wire  fork10_outs_2_valid;
  wire  fork10_outs_2_ready;
  wire [7:0] fork10_outs_3;
  wire  fork10_outs_3_valid;
  wire  fork10_outs_3_ready;
  wire [15:0] extsi14_outs;
  wire  extsi14_outs_valid;
  wire  extsi14_outs_ready;
  wire [15:0] extsi15_outs;
  wire  extsi15_outs_valid;
  wire  extsi15_outs_ready;
  wire [15:0] extsi16_outs;
  wire  extsi16_outs_valid;
  wire  extsi16_outs_ready;
  wire  source0_outs_valid;
  wire  source0_outs_ready;
  wire [1:0] constant2_outs;
  wire  constant2_outs_valid;
  wire  constant2_outs_ready;
  wire [8:0] extui0_outs;
  wire  extui0_outs_valid;
  wire  extui0_outs_ready;
  wire [8:0] addi0_result;
  wire  addi0_result_valid;
  wire  addi0_result_ready;
  wire [8:0] shrsi1_result;
  wire  shrsi1_result_valid;
  wire  shrsi1_result_ready;
  wire [7:0] trunci3_outs;
  wire  trunci3_outs_valid;
  wire  trunci3_outs_ready;
  wire [7:0] fork11_outs_0;
  wire  fork11_outs_0_valid;
  wire  fork11_outs_0_ready;
  wire [7:0] fork11_outs_1;
  wire  fork11_outs_1_valid;
  wire  fork11_outs_1_ready;
  wire [7:0] fork11_outs_2;
  wire  fork11_outs_2_valid;
  wire  fork11_outs_2_ready;
  wire [7:0] fork11_outs_3;
  wire  fork11_outs_3_valid;
  wire  fork11_outs_3_ready;
  wire [15:0] extsi17_outs;
  wire  extsi17_outs_valid;
  wire  extsi17_outs_ready;
  wire [15:0] extsi18_outs;
  wire  extsi18_outs_valid;
  wire  extsi18_outs_ready;
  wire [15:0] muli0_result;
  wire  muli0_result_valid;
  wire  muli0_result_ready;
  wire [15:0] fork12_outs_0;
  wire  fork12_outs_0_valid;
  wire  fork12_outs_0_ready;
  wire [15:0] fork12_outs_1;
  wire  fork12_outs_1_valid;
  wire  fork12_outs_1_ready;
  wire [15:0] fork12_outs_2;
  wire  fork12_outs_2_valid;
  wire  fork12_outs_2_ready;
  wire [0:0] cmpi1_result;
  wire  cmpi1_result_valid;
  wire  cmpi1_result_ready;
  wire [0:0] cmpi2_result;
  wire  cmpi2_result_valid;
  wire  cmpi2_result_ready;
  wire [0:0] fork13_outs_0;
  wire  fork13_outs_0_valid;
  wire  fork13_outs_0_ready;
  wire [0:0] fork13_outs_1;
  wire  fork13_outs_1_valid;
  wire  fork13_outs_1_ready;
  wire [0:0] fork13_outs_2;
  wire  fork13_outs_2_valid;
  wire  fork13_outs_2_ready;
  wire [0:0] fork13_outs_3;
  wire  fork13_outs_3_valid;
  wire  fork13_outs_3_ready;
  wire [0:0] fork13_outs_4;
  wire  fork13_outs_4_valid;
  wire  fork13_outs_4_ready;
  wire [0:0] fork13_outs_5;
  wire  fork13_outs_5_valid;
  wire  fork13_outs_5_ready;
  wire [0:0] fork13_outs_6;
  wire  fork13_outs_6_valid;
  wire  fork13_outs_6_ready;
  wire [0:0] fork13_outs_7;
  wire  fork13_outs_7_valid;
  wire  fork13_outs_7_ready;
  wire [0:0] fork13_outs_8;
  wire  fork13_outs_8_valid;
  wire  fork13_outs_8_ready;
  wire [0:0] fork13_outs_9;
  wire  fork13_outs_9_valid;
  wire  fork13_outs_9_ready;
  wire [0:0] fork13_outs_10;
  wire  fork13_outs_10_valid;
  wire  fork13_outs_10_ready;
  wire [0:0] buffer16_outs;
  wire  buffer16_outs_valid;
  wire  buffer16_outs_ready;
  wire [0:0] buffer17_outs;
  wire  buffer17_outs_valid;
  wire  buffer17_outs_ready;
  wire [0:0] andi1_result;
  wire  andi1_result_valid;
  wire  andi1_result_ready;
  wire [7:0] buffer18_outs;
  wire  buffer18_outs_valid;
  wire  buffer18_outs_ready;
  wire [7:0] buffer19_outs;
  wire  buffer19_outs_valid;
  wire  buffer19_outs_ready;
  wire [7:0] select0_result;
  wire  select0_result_valid;
  wire  select0_result_ready;
  wire [0:0] cmpi3_result;
  wire  cmpi3_result_valid;
  wire  cmpi3_result_ready;
  wire [7:0] cond_br9_trueOut;
  wire  cond_br9_trueOut_valid;
  wire  cond_br9_trueOut_ready;
  wire [7:0] cond_br9_falseOut;
  wire  cond_br9_falseOut_valid;
  wire  cond_br9_falseOut_ready;
  wire [7:0] cond_br10_trueOut;
  wire  cond_br10_trueOut_valid;
  wire  cond_br10_trueOut_ready;
  wire [7:0] cond_br10_falseOut;
  wire  cond_br10_falseOut_valid;
  wire  cond_br10_falseOut_ready;
  wire [7:0] cond_br11_trueOut;
  wire  cond_br11_trueOut_valid;
  wire  cond_br11_trueOut_ready;
  wire [7:0] cond_br11_falseOut;
  wire  cond_br11_falseOut_valid;
  wire  cond_br11_falseOut_ready;
  wire [7:0] cond_br12_trueOut;
  wire  cond_br12_trueOut_valid;
  wire  cond_br12_trueOut_ready;
  wire [7:0] cond_br12_falseOut;
  wire  cond_br12_falseOut_valid;
  wire  cond_br12_falseOut_ready;
  wire [0:0] cond_br13_trueOut;
  wire  cond_br13_trueOut_valid;
  wire  cond_br13_trueOut_ready;
  wire [0:0] cond_br13_falseOut;
  wire  cond_br13_falseOut_valid;
  wire  cond_br13_falseOut_ready;
  wire [0:0] cond_br14_trueOut;
  wire  cond_br14_trueOut_valid;
  wire  cond_br14_trueOut_ready;
  wire [0:0] cond_br14_falseOut;
  wire  cond_br14_falseOut_valid;
  wire  cond_br14_falseOut_ready;
  wire [7:0] cond_br15_trueOut;
  wire  cond_br15_trueOut_valid;
  wire  cond_br15_trueOut_ready;
  wire [7:0] cond_br15_falseOut;
  wire  cond_br15_falseOut_valid;
  wire  cond_br15_falseOut_ready;
  wire [0:0] cond_br16_trueOut;
  wire  cond_br16_trueOut_valid;
  wire  cond_br16_trueOut_ready;
  wire [0:0] cond_br16_falseOut;
  wire  cond_br16_falseOut_valid;
  wire  cond_br16_falseOut_ready;
  wire  buffer24_outs_valid;
  wire  buffer24_outs_ready;
  wire  buffer25_outs_valid;
  wire  buffer25_outs_ready;
  wire  cond_br17_trueOut_valid;
  wire  cond_br17_trueOut_ready;
  wire  cond_br17_falseOut_valid;
  wire  cond_br17_falseOut_ready;
  wire [0:0] buffer40_outs;
  wire  buffer40_outs_valid;
  wire  buffer40_outs_ready;
  wire [0:0] buffer41_outs;
  wire  buffer41_outs_valid;
  wire  buffer41_outs_ready;
  wire [0:0] fork14_outs_0;
  wire  fork14_outs_0_valid;
  wire  fork14_outs_0_ready;
  wire [0:0] fork14_outs_1;
  wire  fork14_outs_1_valid;
  wire  fork14_outs_1_ready;
  wire [0:0] fork14_outs_2;
  wire  fork14_outs_2_valid;
  wire  fork14_outs_2_ready;
  wire [0:0] fork14_outs_3;
  wire  fork14_outs_3_valid;
  wire  fork14_outs_3_ready;
  wire [0:0] fork14_outs_4;
  wire  fork14_outs_4_valid;
  wire  fork14_outs_4_ready;
  wire [0:0] fork14_outs_5;
  wire  fork14_outs_5_valid;
  wire  fork14_outs_5_ready;
  wire [0:0] fork14_outs_6;
  wire  fork14_outs_6_valid;
  wire  fork14_outs_6_ready;
  wire [0:0] fork14_outs_7;
  wire  fork14_outs_7_valid;
  wire  fork14_outs_7_ready;
  wire [7:0] buffer26_outs;
  wire  buffer26_outs_valid;
  wire  buffer26_outs_ready;
  wire [7:0] buffer27_outs;
  wire  buffer27_outs_valid;
  wire  buffer27_outs_ready;
  wire [7:0] cond_br18_trueOut;
  wire  cond_br18_trueOut_valid;
  wire  cond_br18_trueOut_ready;
  wire [7:0] cond_br18_falseOut;
  wire  cond_br18_falseOut_valid;
  wire  cond_br18_falseOut_ready;
  wire [7:0] buffer28_outs;
  wire  buffer28_outs_valid;
  wire  buffer28_outs_ready;
  wire [7:0] buffer29_outs;
  wire  buffer29_outs_valid;
  wire  buffer29_outs_ready;
  wire [7:0] cond_br19_trueOut;
  wire  cond_br19_trueOut_valid;
  wire  cond_br19_trueOut_ready;
  wire [7:0] cond_br19_falseOut;
  wire  cond_br19_falseOut_valid;
  wire  cond_br19_falseOut_ready;
  wire [7:0] buffer32_outs;
  wire  buffer32_outs_valid;
  wire  buffer32_outs_ready;
  wire [7:0] buffer33_outs;
  wire  buffer33_outs_valid;
  wire  buffer33_outs_ready;
  wire [7:0] cond_br20_trueOut;
  wire  cond_br20_trueOut_valid;
  wire  cond_br20_trueOut_ready;
  wire [7:0] cond_br20_falseOut;
  wire  cond_br20_falseOut_valid;
  wire  cond_br20_falseOut_ready;
  wire [0:0] buffer34_outs;
  wire  buffer34_outs_valid;
  wire  buffer34_outs_ready;
  wire [0:0] buffer35_outs;
  wire  buffer35_outs_valid;
  wire  buffer35_outs_ready;
  wire [0:0] cond_br21_trueOut;
  wire  cond_br21_trueOut_valid;
  wire  cond_br21_trueOut_ready;
  wire [0:0] cond_br21_falseOut;
  wire  cond_br21_falseOut_valid;
  wire  cond_br21_falseOut_ready;
  wire [0:0] buffer36_outs;
  wire  buffer36_outs_valid;
  wire  buffer36_outs_ready;
  wire [0:0] buffer37_outs;
  wire  buffer37_outs_valid;
  wire  buffer37_outs_ready;
  wire [0:0] cond_br22_trueOut;
  wire  cond_br22_trueOut_valid;
  wire  cond_br22_trueOut_ready;
  wire [0:0] cond_br22_falseOut;
  wire  cond_br22_falseOut_valid;
  wire  cond_br22_falseOut_ready;
  wire [7:0] buffer38_outs;
  wire  buffer38_outs_valid;
  wire  buffer38_outs_ready;
  wire [7:0] buffer39_outs;
  wire  buffer39_outs_valid;
  wire  buffer39_outs_ready;
  wire [7:0] cond_br23_trueOut;
  wire  cond_br23_trueOut_valid;
  wire  cond_br23_trueOut_ready;
  wire [7:0] cond_br23_falseOut;
  wire  cond_br23_falseOut_valid;
  wire  cond_br23_falseOut_ready;
  wire  buffer42_outs_valid;
  wire  buffer42_outs_ready;
  wire  buffer43_outs_valid;
  wire  buffer43_outs_ready;
  wire  cond_br24_trueOut_valid;
  wire  cond_br24_trueOut_ready;
  wire  cond_br24_falseOut_valid;
  wire  cond_br24_falseOut_ready;
  wire [7:0] buffer30_outs;
  wire  buffer30_outs_valid;
  wire  buffer30_outs_ready;
  wire [7:0] buffer31_outs;
  wire  buffer31_outs_valid;
  wire  buffer31_outs_ready;
  wire [7:0] cond_br25_trueOut;
  wire  cond_br25_trueOut_valid;
  wire  cond_br25_trueOut_ready;
  wire [7:0] cond_br25_falseOut;
  wire  cond_br25_falseOut_valid;
  wire  cond_br25_falseOut_ready;
  wire  source1_outs_valid;
  wire  source1_outs_ready;
  wire [1:0] constant7_outs;
  wire  constant7_outs_valid;
  wire  constant7_outs_ready;
  wire [7:0] extsi19_outs;
  wire  extsi19_outs_valid;
  wire  extsi19_outs_ready;
  wire [7:0] buffer48_outs;
  wire  buffer48_outs_valid;
  wire  buffer48_outs_ready;
  wire [7:0] buffer49_outs;
  wire  buffer49_outs_valid;
  wire  buffer49_outs_ready;
  wire [7:0] addi1_result;
  wire  addi1_result_valid;
  wire  addi1_result_ready;
  wire [7:0] buffer46_outs;
  wire  buffer46_outs_valid;
  wire  buffer46_outs_ready;
  wire [7:0] buffer47_outs;
  wire  buffer47_outs_valid;
  wire  buffer47_outs_ready;
  wire [0:0] buffer52_outs;
  wire  buffer52_outs_valid;
  wire  buffer52_outs_ready;
  wire [0:0] buffer53_outs;
  wire  buffer53_outs_valid;
  wire  buffer53_outs_ready;
  wire [7:0] buffer54_outs;
  wire  buffer54_outs_valid;
  wire  buffer54_outs_ready;
  wire [7:0] buffer55_outs;
  wire  buffer55_outs_valid;
  wire  buffer55_outs_ready;
  wire [0:0] buffer50_outs;
  wire  buffer50_outs_valid;
  wire  buffer50_outs_ready;
  wire [0:0] buffer51_outs;
  wire  buffer51_outs_valid;
  wire  buffer51_outs_ready;
  wire [7:0] buffer44_outs;
  wire  buffer44_outs_valid;
  wire  buffer44_outs_ready;
  wire [7:0] buffer45_outs;
  wire  buffer45_outs_valid;
  wire  buffer45_outs_ready;
  wire  buffer56_outs_valid;
  wire  buffer56_outs_ready;
  wire  buffer57_outs_valid;
  wire  buffer57_outs_ready;
  wire  source2_outs_valid;
  wire  source2_outs_ready;
  wire [31:0] constant6_outs;
  wire  constant6_outs_valid;
  wire  constant6_outs_ready;
  wire [7:0] trunci4_outs;
  wire  trunci4_outs_valid;
  wire  trunci4_outs_ready;
  wire [7:0] buffer62_outs;
  wire  buffer62_outs_valid;
  wire  buffer62_outs_ready;
  wire [7:0] buffer63_outs;
  wire  buffer63_outs_valid;
  wire  buffer63_outs_ready;
  wire [7:0] addi2_result;
  wire  addi2_result_valid;
  wire  addi2_result_ready;
  wire [7:0] buffer60_outs;
  wire  buffer60_outs_valid;
  wire  buffer60_outs_ready;
  wire [7:0] buffer61_outs;
  wire  buffer61_outs_valid;
  wire  buffer61_outs_ready;
  wire [0:0] buffer66_outs;
  wire  buffer66_outs_valid;
  wire  buffer66_outs_ready;
  wire [0:0] buffer67_outs;
  wire  buffer67_outs_valid;
  wire  buffer67_outs_ready;
  wire [7:0] buffer68_outs;
  wire  buffer68_outs_valid;
  wire  buffer68_outs_ready;
  wire [7:0] buffer69_outs;
  wire  buffer69_outs_valid;
  wire  buffer69_outs_ready;
  wire [0:0] buffer64_outs;
  wire  buffer64_outs_valid;
  wire  buffer64_outs_ready;
  wire [0:0] buffer65_outs;
  wire  buffer65_outs_valid;
  wire  buffer65_outs_ready;
  wire [7:0] buffer58_outs;
  wire  buffer58_outs_valid;
  wire  buffer58_outs_ready;
  wire [7:0] buffer59_outs;
  wire  buffer59_outs_valid;
  wire  buffer59_outs_ready;
  wire  buffer70_outs_valid;
  wire  buffer70_outs_ready;
  wire  buffer71_outs_valid;
  wire  buffer71_outs_ready;
  wire [7:0] buffer72_outs;
  wire  buffer72_outs_valid;
  wire  buffer72_outs_ready;
  wire [7:0] buffer73_outs;
  wire  buffer73_outs_valid;
  wire  buffer73_outs_ready;
  wire [0:0] buffer74_outs;
  wire  buffer74_outs_valid;
  wire  buffer74_outs_ready;
  wire [0:0] buffer75_outs;
  wire  buffer75_outs_valid;
  wire  buffer75_outs_ready;
  wire [7:0] buffer76_outs;
  wire  buffer76_outs_valid;
  wire  buffer76_outs_ready;
  wire [7:0] buffer77_outs;
  wire  buffer77_outs_valid;
  wire  buffer77_outs_ready;
  wire [7:0] select1_result;
  wire  select1_result_valid;
  wire  select1_result_ready;

  assign out0 = select1_result;
  assign out0_valid = select1_result_valid;
  assign select1_result_ready = out0_ready;
  assign end_valid = fork0_outs_1_valid;
  assign fork0_outs_1_ready = end_ready;

  fork_dataless #(.SIZE(4)) fork0(
    .ins_valid (start_valid),
    .ins_ready (start_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid ({fork0_outs_3_valid, fork0_outs_2_valid, fork0_outs_1_valid, fork0_outs_0_valid}),
    .outs_ready ({fork0_outs_3_ready, fork0_outs_2_ready, fork0_outs_1_ready, fork0_outs_0_ready})
  );

  fork_type #(.SIZE(2), .DATA_TYPE(8)) fork1(
    .ins (n),
    .ins_valid (n_valid),
    .ins_ready (n_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork1_outs_1, fork1_outs_0}),
    .outs_valid ({fork1_outs_1_valid, fork1_outs_0_valid}),
    .outs_ready ({fork1_outs_1_ready, fork1_outs_0_ready})
  );

  handshake_constant_0 #(.DATA_WIDTH(1)) constant1(
    .ctrl_valid (fork0_outs_0_valid),
    .ctrl_ready (fork0_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant1_outs),
    .outs_valid (constant1_outs_valid),
    .outs_ready (constant1_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(1)) fork2(
    .ins (constant1_outs),
    .ins_valid (constant1_outs_valid),
    .ins_ready (constant1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork2_outs_1, fork2_outs_0}),
    .outs_valid ({fork2_outs_1_valid, fork2_outs_0_valid}),
    .outs_ready ({fork2_outs_1_ready, fork2_outs_0_ready})
  );

  handshake_constant_1 #(.DATA_WIDTH(1)) constant3(
    .ctrl_valid (fork0_outs_3_valid),
    .ctrl_ready (fork0_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant3_outs),
    .outs_valid (constant3_outs_valid),
    .outs_ready (constant3_outs_ready)
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi10(
    .ins (fork2_outs_0),
    .ins_valid (fork2_outs_0_valid),
    .ins_ready (fork2_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi10_outs),
    .outs_valid (extsi10_outs_valid),
    .outs_ready (extsi10_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(1)) fork3(
    .ins (constant3_outs),
    .ins_valid (constant3_outs_valid),
    .ins_ready (constant3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork3_outs_1, fork3_outs_0}),
    .outs_valid ({fork3_outs_1_valid, fork3_outs_0_valid}),
    .outs_ready ({fork3_outs_1_ready, fork3_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(1), .OUTPUT_TYPE(8)) extsi11(
    .ins (fork2_outs_1),
    .ins_valid (fork2_outs_1_valid),
    .ins_ready (fork2_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi11_outs),
    .outs_valid (extsi11_outs_valid),
    .outs_ready (extsi11_outs_ready)
  );

  mux #(.SIZE(4), .DATA_TYPE(8), .SELECT_TYPE(2)) mux0(
    .index (fork6_outs_1),
    .index_valid (fork6_outs_1_valid),
    .index_ready (fork6_outs_1_ready),
    .ins ({addi2_result, buffer47_outs, cond_br10_falseOut, fork1_outs_1}),
    .ins_valid ({addi2_result_valid, buffer47_outs_valid, cond_br10_falseOut_valid, fork1_outs_1_valid}),
    .ins_ready ({addi2_result_ready, buffer47_outs_ready, cond_br10_falseOut_ready, fork1_outs_1_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux0_outs),
    .outs_valid (mux0_outs_valid),
    .outs_ready (mux0_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer0(
    .ins (mux0_outs),
    .ins_valid (mux0_outs_valid),
    .ins_ready (mux0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer0_outs),
    .outs_valid (buffer0_outs_valid),
    .outs_ready (buffer0_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer1(
    .ins (buffer0_outs),
    .ins_valid (buffer0_outs_valid),
    .ins_ready (buffer0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer1_outs),
    .outs_valid (buffer1_outs_valid),
    .outs_ready (buffer1_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(8)) fork4(
    .ins (buffer1_outs),
    .ins_valid (buffer1_outs_valid),
    .ins_ready (buffer1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork4_outs_1, fork4_outs_0}),
    .outs_valid ({fork4_outs_1_valid, fork4_outs_0_valid}),
    .outs_ready ({fork4_outs_1_ready, fork4_outs_0_ready})
  );

  mux #(.SIZE(4), .DATA_TYPE(8), .SELECT_TYPE(2)) mux1(
    .index (fork6_outs_2),
    .index_valid (fork6_outs_2_valid),
    .index_ready (fork6_outs_2_ready),
    .ins ({buffer61_outs, addi1_result, cond_br11_falseOut, extsi10_outs}),
    .ins_valid ({buffer61_outs_valid, addi1_result_valid, cond_br11_falseOut_valid, extsi10_outs_valid}),
    .ins_ready ({buffer61_outs_ready, addi1_result_ready, cond_br11_falseOut_ready, extsi10_outs_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux1_outs),
    .outs_valid (mux1_outs_valid),
    .outs_ready (mux1_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer2(
    .ins (mux1_outs),
    .ins_valid (mux1_outs_valid),
    .ins_ready (mux1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer2_outs),
    .outs_valid (buffer2_outs_valid),
    .outs_ready (buffer2_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer3(
    .ins (buffer2_outs),
    .ins_valid (buffer2_outs_valid),
    .ins_ready (buffer2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer3_outs),
    .outs_valid (buffer3_outs_valid),
    .outs_ready (buffer3_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(8)) fork5(
    .ins (buffer3_outs),
    .ins_valid (buffer3_outs_valid),
    .ins_ready (buffer3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork5_outs_1, fork5_outs_0}),
    .outs_valid ({fork5_outs_1_valid, fork5_outs_0_valid}),
    .outs_ready ({fork5_outs_1_ready, fork5_outs_0_ready})
  );

  mux #(.SIZE(4), .DATA_TYPE(1), .SELECT_TYPE(2)) mux2(
    .index (fork6_outs_3),
    .index_valid (fork6_outs_3_valid),
    .index_ready (fork6_outs_3_ready),
    .ins ({buffer67_outs, buffer53_outs, cond_br14_falseOut, fork3_outs_1}),
    .ins_valid ({buffer67_outs_valid, buffer53_outs_valid, cond_br14_falseOut_valid, fork3_outs_1_valid}),
    .ins_ready ({buffer67_outs_ready, buffer53_outs_ready, cond_br14_falseOut_ready, fork3_outs_1_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux2_outs),
    .outs_valid (mux2_outs_valid),
    .outs_ready (mux2_outs_ready)
  );

  mux #(.SIZE(4), .DATA_TYPE(8), .SELECT_TYPE(2)) mux3(
    .index (fork6_outs_4),
    .index_valid (fork6_outs_4_valid),
    .index_ready (fork6_outs_4_ready),
    .ins ({buffer69_outs, buffer55_outs, cond_br15_falseOut, extsi11_outs}),
    .ins_valid ({buffer69_outs_valid, buffer55_outs_valid, cond_br15_falseOut_valid, extsi11_outs_valid}),
    .ins_ready ({buffer69_outs_ready, buffer55_outs_ready, cond_br15_falseOut_ready, extsi11_outs_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux3_outs),
    .outs_valid (mux3_outs_valid),
    .outs_ready (mux3_outs_ready)
  );

  mux #(.SIZE(4), .DATA_TYPE(1), .SELECT_TYPE(2)) mux4(
    .index (fork6_outs_5),
    .index_valid (fork6_outs_5_valid),
    .index_ready (fork6_outs_5_ready),
    .ins ({buffer65_outs, buffer51_outs, cond_br13_falseOut, fork3_outs_0}),
    .ins_valid ({buffer65_outs_valid, buffer51_outs_valid, cond_br13_falseOut_valid, fork3_outs_0_valid}),
    .ins_ready ({buffer65_outs_ready, buffer51_outs_ready, cond_br13_falseOut_ready, fork3_outs_0_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux4_outs),
    .outs_valid (mux4_outs_valid),
    .outs_ready (mux4_outs_ready)
  );

  mux #(.SIZE(4), .DATA_TYPE(8), .SELECT_TYPE(2)) mux5(
    .index (fork6_outs_0),
    .index_valid (fork6_outs_0_valid),
    .index_ready (fork6_outs_0_ready),
    .ins ({buffer59_outs, buffer45_outs, cond_br9_falseOut, fork1_outs_0}),
    .ins_valid ({buffer59_outs_valid, buffer45_outs_valid, cond_br9_falseOut_valid, fork1_outs_0_valid}),
    .ins_ready ({buffer59_outs_ready, buffer45_outs_ready, cond_br9_falseOut_ready, fork1_outs_0_ready}),
    .clk (clk),
    .rst (rst),
    .outs (mux5_outs),
    .outs_valid (mux5_outs_valid),
    .outs_ready (mux5_outs_ready)
  );

  control_merge_dataless #(.SIZE(4), .INDEX_TYPE(2)) control_merge0(
    .ins_valid ({buffer71_outs_valid, buffer57_outs_valid, cond_br17_falseOut_valid, fork0_outs_2_valid}),
    .ins_ready ({buffer71_outs_ready, buffer57_outs_ready, cond_br17_falseOut_ready, fork0_outs_2_ready}),
    .clk (clk),
    .rst (rst),
    .outs_valid (control_merge0_outs_valid),
    .outs_ready (control_merge0_outs_ready),
    .index (control_merge0_index),
    .index_valid (control_merge0_index_valid),
    .index_ready (control_merge0_index_ready)
  );

  fork_type #(.SIZE(6), .DATA_TYPE(2)) fork6(
    .ins (control_merge0_index),
    .ins_valid (control_merge0_index_valid),
    .ins_ready (control_merge0_index_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork6_outs_5, fork6_outs_4, fork6_outs_3, fork6_outs_2, fork6_outs_1, fork6_outs_0}),
    .outs_valid ({fork6_outs_5_valid, fork6_outs_4_valid, fork6_outs_3_valid, fork6_outs_2_valid, fork6_outs_1_valid, fork6_outs_0_valid}),
    .outs_ready ({fork6_outs_5_ready, fork6_outs_4_ready, fork6_outs_3_ready, fork6_outs_2_ready, fork6_outs_1_ready, fork6_outs_0_ready})
  );

  handshake_cmpi_0 #(.DATA_TYPE(8)) cmpi0(
    .lhs (fork5_outs_0),
    .lhs_valid (fork5_outs_0_valid),
    .lhs_ready (fork5_outs_0_ready),
    .rhs (fork4_outs_0),
    .rhs_valid (fork4_outs_0_valid),
    .rhs_ready (fork4_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi0_result),
    .result_valid (cmpi0_result_valid),
    .result_ready (cmpi0_result_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer8(
    .ins (mux4_outs),
    .ins_valid (mux4_outs_valid),
    .ins_ready (mux4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer8_outs),
    .outs_valid (buffer8_outs_valid),
    .outs_ready (buffer8_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer9(
    .ins (buffer8_outs),
    .ins_valid (buffer8_outs_valid),
    .ins_ready (buffer8_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer9_outs),
    .outs_valid (buffer9_outs_valid),
    .outs_ready (buffer9_outs_ready)
  );

  andi #(.DATA_TYPE(1)) andi0(
    .lhs (cmpi0_result),
    .lhs_valid (cmpi0_result_valid),
    .lhs_ready (cmpi0_result_ready),
    .rhs (buffer9_outs),
    .rhs_valid (buffer9_outs_valid),
    .rhs_ready (buffer9_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (andi0_result),
    .result_valid (andi0_result_valid),
    .result_ready (andi0_result_ready)
  );

  fork_type #(.SIZE(6), .DATA_TYPE(1)) fork7(
    .ins (andi0_result),
    .ins_valid (andi0_result_valid),
    .ins_ready (andi0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork7_outs_5, fork7_outs_4, fork7_outs_3, fork7_outs_2, fork7_outs_1, fork7_outs_0}),
    .outs_valid ({fork7_outs_5_valid, fork7_outs_4_valid, fork7_outs_3_valid, fork7_outs_2_valid, fork7_outs_1_valid, fork7_outs_0_valid}),
    .outs_ready ({fork7_outs_5_ready, fork7_outs_4_ready, fork7_outs_3_ready, fork7_outs_2_ready, fork7_outs_1_ready, fork7_outs_0_ready})
  );

  cond_br #(.DATA_TYPE(8)) cond_br3(
    .condition (fork7_outs_5),
    .condition_valid (fork7_outs_5_valid),
    .condition_ready (fork7_outs_5_ready),
    .data (fork4_outs_1),
    .data_valid (fork4_outs_1_valid),
    .data_ready (fork4_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br3_trueOut),
    .trueOut_valid (cond_br3_trueOut_valid),
    .trueOut_ready (cond_br3_trueOut_ready),
    .falseOut (cond_br3_falseOut),
    .falseOut_valid (cond_br3_falseOut_valid),
    .falseOut_ready (cond_br3_falseOut_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer4(
    .ins (mux2_outs),
    .ins_valid (mux2_outs_valid),
    .ins_ready (mux2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer4_outs),
    .outs_valid (buffer4_outs_valid),
    .outs_ready (buffer4_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer5(
    .ins (buffer4_outs),
    .ins_valid (buffer4_outs_valid),
    .ins_ready (buffer4_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer5_outs),
    .outs_valid (buffer5_outs_valid),
    .outs_ready (buffer5_outs_ready)
  );

  cond_br #(.DATA_TYPE(1)) cond_br4(
    .condition (fork7_outs_4),
    .condition_valid (fork7_outs_4_valid),
    .condition_ready (fork7_outs_4_ready),
    .data (buffer5_outs),
    .data_valid (buffer5_outs_valid),
    .data_ready (buffer5_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br4_trueOut),
    .trueOut_valid (cond_br4_trueOut_valid),
    .trueOut_ready (cond_br4_trueOut_ready),
    .falseOut (cond_br4_falseOut),
    .falseOut_valid (cond_br4_falseOut_valid),
    .falseOut_ready (cond_br4_falseOut_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer6(
    .ins (mux3_outs),
    .ins_valid (mux3_outs_valid),
    .ins_ready (mux3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer6_outs),
    .outs_valid (buffer6_outs_valid),
    .outs_ready (buffer6_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer7(
    .ins (buffer6_outs),
    .ins_valid (buffer6_outs_valid),
    .ins_ready (buffer6_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer7_outs),
    .outs_valid (buffer7_outs_valid),
    .outs_ready (buffer7_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br5(
    .condition (fork7_outs_3),
    .condition_valid (fork7_outs_3_valid),
    .condition_ready (fork7_outs_3_ready),
    .data (buffer7_outs),
    .data_valid (buffer7_outs_valid),
    .data_ready (buffer7_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br5_trueOut),
    .trueOut_valid (cond_br5_trueOut_valid),
    .trueOut_ready (cond_br5_trueOut_ready),
    .falseOut (cond_br5_falseOut),
    .falseOut_valid (cond_br5_falseOut_valid),
    .falseOut_ready (cond_br5_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br6(
    .condition (fork7_outs_2),
    .condition_valid (fork7_outs_2_valid),
    .condition_ready (fork7_outs_2_ready),
    .data (fork5_outs_1),
    .data_valid (fork5_outs_1_valid),
    .data_ready (fork5_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br6_trueOut),
    .trueOut_valid (cond_br6_trueOut_valid),
    .trueOut_ready (cond_br6_trueOut_ready),
    .falseOut (cond_br6_falseOut),
    .falseOut_valid (cond_br6_falseOut_valid),
    .falseOut_ready (cond_br6_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink0(
    .ins (cond_br6_falseOut),
    .ins_valid (cond_br6_falseOut_valid),
    .ins_ready (cond_br6_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(8)) buffer10(
    .ins (mux5_outs),
    .ins_valid (mux5_outs_valid),
    .ins_ready (mux5_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer10_outs),
    .outs_valid (buffer10_outs_valid),
    .outs_ready (buffer10_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer11(
    .ins (buffer10_outs),
    .ins_valid (buffer10_outs_valid),
    .ins_ready (buffer10_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer11_outs),
    .outs_valid (buffer11_outs_valid),
    .outs_ready (buffer11_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br7(
    .condition (fork7_outs_0),
    .condition_valid (fork7_outs_0_valid),
    .condition_ready (fork7_outs_0_ready),
    .data (buffer11_outs),
    .data_valid (buffer11_outs_valid),
    .data_ready (buffer11_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br7_trueOut),
    .trueOut_valid (cond_br7_trueOut_valid),
    .trueOut_ready (cond_br7_trueOut_ready),
    .falseOut (cond_br7_falseOut),
    .falseOut_valid (cond_br7_falseOut_valid),
    .falseOut_ready (cond_br7_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink1(
    .ins (cond_br7_falseOut),
    .ins_valid (cond_br7_falseOut_valid),
    .ins_ready (cond_br7_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb_dataless buffer12(
    .ins_valid (control_merge0_outs_valid),
    .ins_ready (control_merge0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer12_outs_valid),
    .outs_ready (buffer12_outs_ready)
  );

  tehb_dataless buffer13(
    .ins_valid (buffer12_outs_valid),
    .ins_ready (buffer12_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer13_outs_valid),
    .outs_ready (buffer13_outs_ready)
  );

  cond_br_dataless cond_br8(
    .condition (fork7_outs_1),
    .condition_valid (fork7_outs_1_valid),
    .condition_ready (fork7_outs_1_ready),
    .data_valid (buffer13_outs_valid),
    .data_ready (buffer13_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br8_trueOut_valid),
    .trueOut_ready (cond_br8_trueOut_ready),
    .falseOut_valid (cond_br8_falseOut_valid),
    .falseOut_ready (cond_br8_falseOut_ready)
  );

  sink_dataless sink2(
    .ins_valid (cond_br8_falseOut_valid),
    .ins_ready (cond_br8_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(8)) buffer14(
    .ins (cond_br3_trueOut),
    .ins_valid (cond_br3_trueOut_valid),
    .ins_ready (cond_br3_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer14_outs),
    .outs_valid (buffer14_outs_valid),
    .outs_ready (buffer14_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer15(
    .ins (buffer14_outs),
    .ins_valid (buffer14_outs_valid),
    .ins_ready (buffer14_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer15_outs),
    .outs_valid (buffer15_outs_valid),
    .outs_ready (buffer15_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(8)) fork8(
    .ins (buffer15_outs),
    .ins_valid (buffer15_outs_valid),
    .ins_ready (buffer15_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork8_outs_1, fork8_outs_0}),
    .outs_valid ({fork8_outs_1_valid, fork8_outs_0_valid}),
    .outs_ready ({fork8_outs_1_ready, fork8_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(9)) extsi12(
    .ins (fork8_outs_0),
    .ins_valid (fork8_outs_0_valid),
    .ins_ready (fork8_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi12_outs),
    .outs_valid (extsi12_outs_valid),
    .outs_ready (extsi12_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer20(
    .ins (cond_br6_trueOut),
    .ins_valid (cond_br6_trueOut_valid),
    .ins_ready (cond_br6_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer20_outs),
    .outs_valid (buffer20_outs_valid),
    .outs_ready (buffer20_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer21(
    .ins (buffer20_outs),
    .ins_valid (buffer20_outs_valid),
    .ins_ready (buffer20_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer21_outs),
    .outs_valid (buffer21_outs_valid),
    .outs_ready (buffer21_outs_ready)
  );

  fork_type #(.SIZE(2), .DATA_TYPE(8)) fork9(
    .ins (buffer21_outs),
    .ins_valid (buffer21_outs_valid),
    .ins_ready (buffer21_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork9_outs_1, fork9_outs_0}),
    .outs_valid ({fork9_outs_1_valid, fork9_outs_0_valid}),
    .outs_ready ({fork9_outs_1_ready, fork9_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(9)) extsi13(
    .ins (fork9_outs_0),
    .ins_valid (fork9_outs_0_valid),
    .ins_ready (fork9_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi13_outs),
    .outs_valid (extsi13_outs_valid),
    .outs_ready (extsi13_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer22(
    .ins (cond_br7_trueOut),
    .ins_valid (cond_br7_trueOut_valid),
    .ins_ready (cond_br7_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer22_outs),
    .outs_valid (buffer22_outs_valid),
    .outs_ready (buffer22_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer23(
    .ins (buffer22_outs),
    .ins_valid (buffer22_outs_valid),
    .ins_ready (buffer22_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer23_outs),
    .outs_valid (buffer23_outs_valid),
    .outs_ready (buffer23_outs_ready)
  );

  fork_type #(.SIZE(4), .DATA_TYPE(8)) fork10(
    .ins (buffer23_outs),
    .ins_valid (buffer23_outs_valid),
    .ins_ready (buffer23_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork10_outs_3, fork10_outs_2, fork10_outs_1, fork10_outs_0}),
    .outs_valid ({fork10_outs_3_valid, fork10_outs_2_valid, fork10_outs_1_valid, fork10_outs_0_valid}),
    .outs_ready ({fork10_outs_3_ready, fork10_outs_2_ready, fork10_outs_1_ready, fork10_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(16)) extsi14(
    .ins (fork10_outs_1),
    .ins_valid (fork10_outs_1_valid),
    .ins_ready (fork10_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi14_outs),
    .outs_valid (extsi14_outs_valid),
    .outs_ready (extsi14_outs_ready)
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(16)) extsi15(
    .ins (fork10_outs_2),
    .ins_valid (fork10_outs_2_valid),
    .ins_ready (fork10_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi15_outs),
    .outs_valid (extsi15_outs_valid),
    .outs_ready (extsi15_outs_ready)
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(16)) extsi16(
    .ins (fork10_outs_3),
    .ins_valid (fork10_outs_3_valid),
    .ins_ready (fork10_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi16_outs),
    .outs_valid (extsi16_outs_valid),
    .outs_ready (extsi16_outs_ready)
  );

  source source0(
    .clk (clk),
    .rst (rst),
    .outs_valid (source0_outs_valid),
    .outs_ready (source0_outs_ready)
  );

  handshake_constant_2 #(.DATA_WIDTH(2)) constant2(
    .ctrl_valid (source0_outs_valid),
    .ctrl_ready (source0_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant2_outs),
    .outs_valid (constant2_outs_valid),
    .outs_ready (constant2_outs_ready)
  );

  extui #(.INPUT_TYPE(2), .OUTPUT_TYPE(9)) extui0(
    .ins (constant2_outs),
    .ins_valid (constant2_outs_valid),
    .ins_ready (constant2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extui0_outs),
    .outs_valid (extui0_outs_valid),
    .outs_ready (extui0_outs_ready)
  );

  addi #(.DATA_TYPE(9)) addi0(
    .lhs (extsi13_outs),
    .lhs_valid (extsi13_outs_valid),
    .lhs_ready (extsi13_outs_ready),
    .rhs (extsi12_outs),
    .rhs_valid (extsi12_outs_valid),
    .rhs_ready (extsi12_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi0_result),
    .result_valid (addi0_result_valid),
    .result_ready (addi0_result_ready)
  );

  shrsi #(.DATA_TYPE(9)) shrsi1(
    .lhs (addi0_result),
    .lhs_valid (addi0_result_valid),
    .lhs_ready (addi0_result_ready),
    .rhs (extui0_outs),
    .rhs_valid (extui0_outs_valid),
    .rhs_ready (extui0_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (shrsi1_result),
    .result_valid (shrsi1_result_valid),
    .result_ready (shrsi1_result_ready)
  );

  trunci #(.INPUT_TYPE(9), .OUTPUT_TYPE(8)) trunci3(
    .ins (shrsi1_result),
    .ins_valid (shrsi1_result_valid),
    .ins_ready (shrsi1_result_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci3_outs),
    .outs_valid (trunci3_outs_valid),
    .outs_ready (trunci3_outs_ready)
  );

  fork_type #(.SIZE(4), .DATA_TYPE(8)) fork11(
    .ins (trunci3_outs),
    .ins_valid (trunci3_outs_valid),
    .ins_ready (trunci3_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork11_outs_3, fork11_outs_2, fork11_outs_1, fork11_outs_0}),
    .outs_valid ({fork11_outs_3_valid, fork11_outs_2_valid, fork11_outs_1_valid, fork11_outs_0_valid}),
    .outs_ready ({fork11_outs_3_ready, fork11_outs_2_ready, fork11_outs_1_ready, fork11_outs_0_ready})
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(16)) extsi17(
    .ins (fork11_outs_3),
    .ins_valid (fork11_outs_3_valid),
    .ins_ready (fork11_outs_3_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi17_outs),
    .outs_valid (extsi17_outs_valid),
    .outs_ready (extsi17_outs_ready)
  );

  extsi #(.INPUT_TYPE(8), .OUTPUT_TYPE(16)) extsi18(
    .ins (fork11_outs_2),
    .ins_valid (fork11_outs_2_valid),
    .ins_ready (fork11_outs_2_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi18_outs),
    .outs_valid (extsi18_outs_valid),
    .outs_ready (extsi18_outs_ready)
  );

  muli #(.DATA_TYPE(16)) muli0(
    .lhs (extsi18_outs),
    .lhs_valid (extsi18_outs_valid),
    .lhs_ready (extsi18_outs_ready),
    .rhs (extsi17_outs),
    .rhs_valid (extsi17_outs_valid),
    .rhs_ready (extsi17_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (muli0_result),
    .result_valid (muli0_result_valid),
    .result_ready (muli0_result_ready)
  );

  fork_type #(.SIZE(3), .DATA_TYPE(16)) fork12(
    .ins (muli0_result),
    .ins_valid (muli0_result_valid),
    .ins_ready (muli0_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork12_outs_2, fork12_outs_1, fork12_outs_0}),
    .outs_valid ({fork12_outs_2_valid, fork12_outs_1_valid, fork12_outs_0_valid}),
    .outs_ready ({fork12_outs_2_ready, fork12_outs_1_ready, fork12_outs_0_ready})
  );

  handshake_cmpi_1 #(.DATA_TYPE(16)) cmpi1(
    .lhs (fork12_outs_2),
    .lhs_valid (fork12_outs_2_valid),
    .lhs_ready (fork12_outs_2_ready),
    .rhs (extsi16_outs),
    .rhs_valid (extsi16_outs_valid),
    .rhs_ready (extsi16_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi1_result),
    .result_valid (cmpi1_result_valid),
    .result_ready (cmpi1_result_ready)
  );

  handshake_cmpi_2 #(.DATA_TYPE(16)) cmpi2(
    .lhs (fork12_outs_1),
    .lhs_valid (fork12_outs_1_valid),
    .lhs_ready (fork12_outs_1_ready),
    .rhs (extsi15_outs),
    .rhs_valid (extsi15_outs_valid),
    .rhs_ready (extsi15_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi2_result),
    .result_valid (cmpi2_result_valid),
    .result_ready (cmpi2_result_ready)
  );

  fork_type #(.SIZE(11), .DATA_TYPE(1)) fork13(
    .ins (cmpi2_result),
    .ins_valid (cmpi2_result_valid),
    .ins_ready (cmpi2_result_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork13_outs_10, fork13_outs_9, fork13_outs_8, fork13_outs_7, fork13_outs_6, fork13_outs_5, fork13_outs_4, fork13_outs_3, fork13_outs_2, fork13_outs_1, fork13_outs_0}),
    .outs_valid ({fork13_outs_10_valid, fork13_outs_9_valid, fork13_outs_8_valid, fork13_outs_7_valid, fork13_outs_6_valid, fork13_outs_5_valid, fork13_outs_4_valid, fork13_outs_3_valid, fork13_outs_2_valid, fork13_outs_1_valid, fork13_outs_0_valid}),
    .outs_ready ({fork13_outs_10_ready, fork13_outs_9_ready, fork13_outs_8_ready, fork13_outs_7_ready, fork13_outs_6_ready, fork13_outs_5_ready, fork13_outs_4_ready, fork13_outs_3_ready, fork13_outs_2_ready, fork13_outs_1_ready, fork13_outs_0_ready})
  );

  oehb #(.DATA_TYPE(1)) buffer16(
    .ins (cond_br4_trueOut),
    .ins_valid (cond_br4_trueOut_valid),
    .ins_ready (cond_br4_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer16_outs),
    .outs_valid (buffer16_outs_valid),
    .outs_ready (buffer16_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer17(
    .ins (buffer16_outs),
    .ins_valid (buffer16_outs_valid),
    .ins_ready (buffer16_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer17_outs),
    .outs_valid (buffer17_outs_valid),
    .outs_ready (buffer17_outs_ready)
  );

  andi #(.DATA_TYPE(1)) andi1(
    .lhs (fork13_outs_1),
    .lhs_valid (fork13_outs_1_valid),
    .lhs_ready (fork13_outs_1_ready),
    .rhs (buffer17_outs),
    .rhs_valid (buffer17_outs_valid),
    .rhs_ready (buffer17_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (andi1_result),
    .result_valid (andi1_result_valid),
    .result_ready (andi1_result_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer18(
    .ins (cond_br5_trueOut),
    .ins_valid (cond_br5_trueOut_valid),
    .ins_ready (cond_br5_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer18_outs),
    .outs_valid (buffer18_outs_valid),
    .outs_ready (buffer18_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer19(
    .ins (buffer18_outs),
    .ins_valid (buffer18_outs_valid),
    .ins_ready (buffer18_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer19_outs),
    .outs_valid (buffer19_outs_valid),
    .outs_ready (buffer19_outs_ready)
  );

  selector #(.DATA_TYPE(8)) select0(
    .condition (cmpi1_result),
    .condition_valid (cmpi1_result_valid),
    .condition_ready (cmpi1_result_ready),
    .trueValue (fork11_outs_0),
    .trueValue_valid (fork11_outs_0_valid),
    .trueValue_ready (fork11_outs_0_ready),
    .falseValue (buffer19_outs),
    .falseValue_valid (buffer19_outs_valid),
    .falseValue_ready (buffer19_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (select0_result),
    .result_valid (select0_result_valid),
    .result_ready (select0_result_ready)
  );

  handshake_cmpi_3 #(.DATA_TYPE(16)) cmpi3(
    .lhs (fork12_outs_0),
    .lhs_valid (fork12_outs_0_valid),
    .lhs_ready (fork12_outs_0_ready),
    .rhs (extsi14_outs),
    .rhs_valid (extsi14_outs_valid),
    .rhs_ready (extsi14_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (cmpi3_result),
    .result_valid (cmpi3_result_valid),
    .result_ready (cmpi3_result_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br9(
    .condition (fork13_outs_0),
    .condition_valid (fork13_outs_0_valid),
    .condition_ready (fork13_outs_0_ready),
    .data (fork10_outs_0),
    .data_valid (fork10_outs_0_valid),
    .data_ready (fork10_outs_0_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br9_trueOut),
    .trueOut_valid (cond_br9_trueOut_valid),
    .trueOut_ready (cond_br9_trueOut_ready),
    .falseOut (cond_br9_falseOut),
    .falseOut_valid (cond_br9_falseOut_valid),
    .falseOut_ready (cond_br9_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br10(
    .condition (fork13_outs_2),
    .condition_valid (fork13_outs_2_valid),
    .condition_ready (fork13_outs_2_ready),
    .data (fork8_outs_1),
    .data_valid (fork8_outs_1_valid),
    .data_ready (fork8_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br10_trueOut),
    .trueOut_valid (cond_br10_trueOut_valid),
    .trueOut_ready (cond_br10_trueOut_ready),
    .falseOut (cond_br10_falseOut),
    .falseOut_valid (cond_br10_falseOut_valid),
    .falseOut_ready (cond_br10_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br11(
    .condition (fork13_outs_3),
    .condition_valid (fork13_outs_3_valid),
    .condition_ready (fork13_outs_3_ready),
    .data (fork9_outs_1),
    .data_valid (fork9_outs_1_valid),
    .data_ready (fork9_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br11_trueOut),
    .trueOut_valid (cond_br11_trueOut_valid),
    .trueOut_ready (cond_br11_trueOut_ready),
    .falseOut (cond_br11_falseOut),
    .falseOut_valid (cond_br11_falseOut_valid),
    .falseOut_ready (cond_br11_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br12(
    .condition (fork13_outs_10),
    .condition_valid (fork13_outs_10_valid),
    .condition_ready (fork13_outs_10_ready),
    .data (fork11_outs_1),
    .data_valid (fork11_outs_1_valid),
    .data_ready (fork11_outs_1_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br12_trueOut),
    .trueOut_valid (cond_br12_trueOut_valid),
    .trueOut_ready (cond_br12_trueOut_ready),
    .falseOut (cond_br12_falseOut),
    .falseOut_valid (cond_br12_falseOut_valid),
    .falseOut_ready (cond_br12_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink4(
    .ins (cond_br12_falseOut),
    .ins_valid (cond_br12_falseOut_valid),
    .ins_ready (cond_br12_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  cond_br #(.DATA_TYPE(1)) cond_br13(
    .condition (fork13_outs_4),
    .condition_valid (fork13_outs_4_valid),
    .condition_ready (fork13_outs_4_ready),
    .data (fork13_outs_5),
    .data_valid (fork13_outs_5_valid),
    .data_ready (fork13_outs_5_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br13_trueOut),
    .trueOut_valid (cond_br13_trueOut_valid),
    .trueOut_ready (cond_br13_trueOut_ready),
    .falseOut (cond_br13_falseOut),
    .falseOut_valid (cond_br13_falseOut_valid),
    .falseOut_ready (cond_br13_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(1)) cond_br14(
    .condition (fork13_outs_6),
    .condition_valid (fork13_outs_6_valid),
    .condition_ready (fork13_outs_6_ready),
    .data (andi1_result),
    .data_valid (andi1_result_valid),
    .data_ready (andi1_result_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br14_trueOut),
    .trueOut_valid (cond_br14_trueOut_valid),
    .trueOut_ready (cond_br14_trueOut_ready),
    .falseOut (cond_br14_falseOut),
    .falseOut_valid (cond_br14_falseOut_valid),
    .falseOut_ready (cond_br14_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br15(
    .condition (fork13_outs_7),
    .condition_valid (fork13_outs_7_valid),
    .condition_ready (fork13_outs_7_ready),
    .data (select0_result),
    .data_valid (select0_result_valid),
    .data_ready (select0_result_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br15_trueOut),
    .trueOut_valid (cond_br15_trueOut_valid),
    .trueOut_ready (cond_br15_trueOut_ready),
    .falseOut (cond_br15_falseOut),
    .falseOut_valid (cond_br15_falseOut_valid),
    .falseOut_ready (cond_br15_falseOut_ready)
  );

  cond_br #(.DATA_TYPE(1)) cond_br16(
    .condition (fork13_outs_8),
    .condition_valid (fork13_outs_8_valid),
    .condition_ready (fork13_outs_8_ready),
    .data (cmpi3_result),
    .data_valid (cmpi3_result_valid),
    .data_ready (cmpi3_result_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br16_trueOut),
    .trueOut_valid (cond_br16_trueOut_valid),
    .trueOut_ready (cond_br16_trueOut_ready),
    .falseOut (cond_br16_falseOut),
    .falseOut_valid (cond_br16_falseOut_valid),
    .falseOut_ready (cond_br16_falseOut_ready)
  );

  sink #(.DATA_TYPE(1)) sink5(
    .ins (cond_br16_falseOut),
    .ins_valid (cond_br16_falseOut_valid),
    .ins_ready (cond_br16_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb_dataless buffer24(
    .ins_valid (cond_br8_trueOut_valid),
    .ins_ready (cond_br8_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer24_outs_valid),
    .outs_ready (buffer24_outs_ready)
  );

  tehb_dataless buffer25(
    .ins_valid (buffer24_outs_valid),
    .ins_ready (buffer24_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer25_outs_valid),
    .outs_ready (buffer25_outs_ready)
  );

  cond_br_dataless cond_br17(
    .condition (fork13_outs_9),
    .condition_valid (fork13_outs_9_valid),
    .condition_ready (fork13_outs_9_ready),
    .data_valid (buffer25_outs_valid),
    .data_ready (buffer25_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br17_trueOut_valid),
    .trueOut_ready (cond_br17_trueOut_ready),
    .falseOut_valid (cond_br17_falseOut_valid),
    .falseOut_ready (cond_br17_falseOut_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer40(
    .ins (cond_br16_trueOut),
    .ins_valid (cond_br16_trueOut_valid),
    .ins_ready (cond_br16_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer40_outs),
    .outs_valid (buffer40_outs_valid),
    .outs_ready (buffer40_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer41(
    .ins (buffer40_outs),
    .ins_valid (buffer40_outs_valid),
    .ins_ready (buffer40_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer41_outs),
    .outs_valid (buffer41_outs_valid),
    .outs_ready (buffer41_outs_ready)
  );

  fork_type #(.SIZE(8), .DATA_TYPE(1)) fork14(
    .ins (buffer41_outs),
    .ins_valid (buffer41_outs_valid),
    .ins_ready (buffer41_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs ({fork14_outs_7, fork14_outs_6, fork14_outs_5, fork14_outs_4, fork14_outs_3, fork14_outs_2, fork14_outs_1, fork14_outs_0}),
    .outs_valid ({fork14_outs_7_valid, fork14_outs_6_valid, fork14_outs_5_valid, fork14_outs_4_valid, fork14_outs_3_valid, fork14_outs_2_valid, fork14_outs_1_valid, fork14_outs_0_valid}),
    .outs_ready ({fork14_outs_7_ready, fork14_outs_6_ready, fork14_outs_5_ready, fork14_outs_4_ready, fork14_outs_3_ready, fork14_outs_2_ready, fork14_outs_1_ready, fork14_outs_0_ready})
  );

  oehb #(.DATA_TYPE(8)) buffer26(
    .ins (cond_br9_trueOut),
    .ins_valid (cond_br9_trueOut_valid),
    .ins_ready (cond_br9_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer26_outs),
    .outs_valid (buffer26_outs_valid),
    .outs_ready (buffer26_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer27(
    .ins (buffer26_outs),
    .ins_valid (buffer26_outs_valid),
    .ins_ready (buffer26_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer27_outs),
    .outs_valid (buffer27_outs_valid),
    .outs_ready (buffer27_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br18(
    .condition (fork14_outs_0),
    .condition_valid (fork14_outs_0_valid),
    .condition_ready (fork14_outs_0_ready),
    .data (buffer27_outs),
    .data_valid (buffer27_outs_valid),
    .data_ready (buffer27_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br18_trueOut),
    .trueOut_valid (cond_br18_trueOut_valid),
    .trueOut_ready (cond_br18_trueOut_ready),
    .falseOut (cond_br18_falseOut),
    .falseOut_valid (cond_br18_falseOut_valid),
    .falseOut_ready (cond_br18_falseOut_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer28(
    .ins (cond_br10_trueOut),
    .ins_valid (cond_br10_trueOut_valid),
    .ins_ready (cond_br10_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer28_outs),
    .outs_valid (buffer28_outs_valid),
    .outs_ready (buffer28_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer29(
    .ins (buffer28_outs),
    .ins_valid (buffer28_outs_valid),
    .ins_ready (buffer28_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer29_outs),
    .outs_valid (buffer29_outs_valid),
    .outs_ready (buffer29_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br19(
    .condition (fork14_outs_7),
    .condition_valid (fork14_outs_7_valid),
    .condition_ready (fork14_outs_7_ready),
    .data (buffer29_outs),
    .data_valid (buffer29_outs_valid),
    .data_ready (buffer29_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br19_trueOut),
    .trueOut_valid (cond_br19_trueOut_valid),
    .trueOut_ready (cond_br19_trueOut_ready),
    .falseOut (cond_br19_falseOut),
    .falseOut_valid (cond_br19_falseOut_valid),
    .falseOut_ready (cond_br19_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink7(
    .ins (cond_br19_falseOut),
    .ins_valid (cond_br19_falseOut_valid),
    .ins_ready (cond_br19_falseOut_ready),
    .clk (clk),
    .rst (rst)
  );

  oehb #(.DATA_TYPE(8)) buffer32(
    .ins (cond_br12_trueOut),
    .ins_valid (cond_br12_trueOut_valid),
    .ins_ready (cond_br12_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer32_outs),
    .outs_valid (buffer32_outs_valid),
    .outs_ready (buffer32_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer33(
    .ins (buffer32_outs),
    .ins_valid (buffer32_outs_valid),
    .ins_ready (buffer32_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer33_outs),
    .outs_valid (buffer33_outs_valid),
    .outs_ready (buffer33_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br20(
    .condition (fork14_outs_1),
    .condition_valid (fork14_outs_1_valid),
    .condition_ready (fork14_outs_1_ready),
    .data (buffer33_outs),
    .data_valid (buffer33_outs_valid),
    .data_ready (buffer33_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br20_trueOut),
    .trueOut_valid (cond_br20_trueOut_valid),
    .trueOut_ready (cond_br20_trueOut_ready),
    .falseOut (cond_br20_falseOut),
    .falseOut_valid (cond_br20_falseOut_valid),
    .falseOut_ready (cond_br20_falseOut_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer34(
    .ins (cond_br13_trueOut),
    .ins_valid (cond_br13_trueOut_valid),
    .ins_ready (cond_br13_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer34_outs),
    .outs_valid (buffer34_outs_valid),
    .outs_ready (buffer34_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer35(
    .ins (buffer34_outs),
    .ins_valid (buffer34_outs_valid),
    .ins_ready (buffer34_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer35_outs),
    .outs_valid (buffer35_outs_valid),
    .outs_ready (buffer35_outs_ready)
  );

  cond_br #(.DATA_TYPE(1)) cond_br21(
    .condition (fork14_outs_6),
    .condition_valid (fork14_outs_6_valid),
    .condition_ready (fork14_outs_6_ready),
    .data (buffer35_outs),
    .data_valid (buffer35_outs_valid),
    .data_ready (buffer35_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br21_trueOut),
    .trueOut_valid (cond_br21_trueOut_valid),
    .trueOut_ready (cond_br21_trueOut_ready),
    .falseOut (cond_br21_falseOut),
    .falseOut_valid (cond_br21_falseOut_valid),
    .falseOut_ready (cond_br21_falseOut_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer36(
    .ins (cond_br14_trueOut),
    .ins_valid (cond_br14_trueOut_valid),
    .ins_ready (cond_br14_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer36_outs),
    .outs_valid (buffer36_outs_valid),
    .outs_ready (buffer36_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer37(
    .ins (buffer36_outs),
    .ins_valid (buffer36_outs_valid),
    .ins_ready (buffer36_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer37_outs),
    .outs_valid (buffer37_outs_valid),
    .outs_ready (buffer37_outs_ready)
  );

  cond_br #(.DATA_TYPE(1)) cond_br22(
    .condition (fork14_outs_5),
    .condition_valid (fork14_outs_5_valid),
    .condition_ready (fork14_outs_5_ready),
    .data (buffer37_outs),
    .data_valid (buffer37_outs_valid),
    .data_ready (buffer37_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br22_trueOut),
    .trueOut_valid (cond_br22_trueOut_valid),
    .trueOut_ready (cond_br22_trueOut_ready),
    .falseOut (cond_br22_falseOut),
    .falseOut_valid (cond_br22_falseOut_valid),
    .falseOut_ready (cond_br22_falseOut_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer38(
    .ins (cond_br15_trueOut),
    .ins_valid (cond_br15_trueOut_valid),
    .ins_ready (cond_br15_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer38_outs),
    .outs_valid (buffer38_outs_valid),
    .outs_ready (buffer38_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer39(
    .ins (buffer38_outs),
    .ins_valid (buffer38_outs_valid),
    .ins_ready (buffer38_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer39_outs),
    .outs_valid (buffer39_outs_valid),
    .outs_ready (buffer39_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br23(
    .condition (fork14_outs_4),
    .condition_valid (fork14_outs_4_valid),
    .condition_ready (fork14_outs_4_ready),
    .data (buffer39_outs),
    .data_valid (buffer39_outs_valid),
    .data_ready (buffer39_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br23_trueOut),
    .trueOut_valid (cond_br23_trueOut_valid),
    .trueOut_ready (cond_br23_trueOut_ready),
    .falseOut (cond_br23_falseOut),
    .falseOut_valid (cond_br23_falseOut_valid),
    .falseOut_ready (cond_br23_falseOut_ready)
  );

  oehb_dataless buffer42(
    .ins_valid (cond_br17_trueOut_valid),
    .ins_ready (cond_br17_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer42_outs_valid),
    .outs_ready (buffer42_outs_ready)
  );

  tehb_dataless buffer43(
    .ins_valid (buffer42_outs_valid),
    .ins_ready (buffer42_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer43_outs_valid),
    .outs_ready (buffer43_outs_ready)
  );

  cond_br_dataless cond_br24(
    .condition (fork14_outs_3),
    .condition_valid (fork14_outs_3_valid),
    .condition_ready (fork14_outs_3_ready),
    .data_valid (buffer43_outs_valid),
    .data_ready (buffer43_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut_valid (cond_br24_trueOut_valid),
    .trueOut_ready (cond_br24_trueOut_ready),
    .falseOut_valid (cond_br24_falseOut_valid),
    .falseOut_ready (cond_br24_falseOut_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer30(
    .ins (cond_br11_trueOut),
    .ins_valid (cond_br11_trueOut_valid),
    .ins_ready (cond_br11_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer30_outs),
    .outs_valid (buffer30_outs_valid),
    .outs_ready (buffer30_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer31(
    .ins (buffer30_outs),
    .ins_valid (buffer30_outs_valid),
    .ins_ready (buffer30_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer31_outs),
    .outs_valid (buffer31_outs_valid),
    .outs_ready (buffer31_outs_ready)
  );

  cond_br #(.DATA_TYPE(8)) cond_br25(
    .condition (fork14_outs_2),
    .condition_valid (fork14_outs_2_valid),
    .condition_ready (fork14_outs_2_ready),
    .data (buffer31_outs),
    .data_valid (buffer31_outs_valid),
    .data_ready (buffer31_outs_ready),
    .clk (clk),
    .rst (rst),
    .trueOut (cond_br25_trueOut),
    .trueOut_valid (cond_br25_trueOut_valid),
    .trueOut_ready (cond_br25_trueOut_ready),
    .falseOut (cond_br25_falseOut),
    .falseOut_valid (cond_br25_falseOut_valid),
    .falseOut_ready (cond_br25_falseOut_ready)
  );

  sink #(.DATA_TYPE(8)) sink8(
    .ins (cond_br25_trueOut),
    .ins_valid (cond_br25_trueOut_valid),
    .ins_ready (cond_br25_trueOut_ready),
    .clk (clk),
    .rst (rst)
  );

  source source1(
    .clk (clk),
    .rst (rst),
    .outs_valid (source1_outs_valid),
    .outs_ready (source1_outs_ready)
  );

  handshake_constant_2 #(.DATA_WIDTH(2)) constant7(
    .ctrl_valid (source1_outs_valid),
    .ctrl_ready (source1_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant7_outs),
    .outs_valid (constant7_outs_valid),
    .outs_ready (constant7_outs_ready)
  );

  extsi #(.INPUT_TYPE(2), .OUTPUT_TYPE(8)) extsi19(
    .ins (constant7_outs),
    .ins_valid (constant7_outs_valid),
    .ins_ready (constant7_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (extsi19_outs),
    .outs_valid (extsi19_outs_valid),
    .outs_ready (extsi19_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer48(
    .ins (cond_br20_trueOut),
    .ins_valid (cond_br20_trueOut_valid),
    .ins_ready (cond_br20_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer48_outs),
    .outs_valid (buffer48_outs_valid),
    .outs_ready (buffer48_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer49(
    .ins (buffer48_outs),
    .ins_valid (buffer48_outs_valid),
    .ins_ready (buffer48_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer49_outs),
    .outs_valid (buffer49_outs_valid),
    .outs_ready (buffer49_outs_ready)
  );

  addi #(.DATA_TYPE(8)) addi1(
    .lhs (buffer49_outs),
    .lhs_valid (buffer49_outs_valid),
    .lhs_ready (buffer49_outs_ready),
    .rhs (extsi19_outs),
    .rhs_valid (extsi19_outs_valid),
    .rhs_ready (extsi19_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi1_result),
    .result_valid (addi1_result_valid),
    .result_ready (addi1_result_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer46(
    .ins (cond_br19_trueOut),
    .ins_valid (cond_br19_trueOut_valid),
    .ins_ready (cond_br19_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer46_outs),
    .outs_valid (buffer46_outs_valid),
    .outs_ready (buffer46_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer47(
    .ins (buffer46_outs),
    .ins_valid (buffer46_outs_valid),
    .ins_ready (buffer46_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer47_outs),
    .outs_valid (buffer47_outs_valid),
    .outs_ready (buffer47_outs_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer52(
    .ins (cond_br22_trueOut),
    .ins_valid (cond_br22_trueOut_valid),
    .ins_ready (cond_br22_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer52_outs),
    .outs_valid (buffer52_outs_valid),
    .outs_ready (buffer52_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer53(
    .ins (buffer52_outs),
    .ins_valid (buffer52_outs_valid),
    .ins_ready (buffer52_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer53_outs),
    .outs_valid (buffer53_outs_valid),
    .outs_ready (buffer53_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer54(
    .ins (cond_br23_trueOut),
    .ins_valid (cond_br23_trueOut_valid),
    .ins_ready (cond_br23_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer54_outs),
    .outs_valid (buffer54_outs_valid),
    .outs_ready (buffer54_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer55(
    .ins (buffer54_outs),
    .ins_valid (buffer54_outs_valid),
    .ins_ready (buffer54_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer55_outs),
    .outs_valid (buffer55_outs_valid),
    .outs_ready (buffer55_outs_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer50(
    .ins (cond_br21_trueOut),
    .ins_valid (cond_br21_trueOut_valid),
    .ins_ready (cond_br21_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer50_outs),
    .outs_valid (buffer50_outs_valid),
    .outs_ready (buffer50_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer51(
    .ins (buffer50_outs),
    .ins_valid (buffer50_outs_valid),
    .ins_ready (buffer50_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer51_outs),
    .outs_valid (buffer51_outs_valid),
    .outs_ready (buffer51_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer44(
    .ins (cond_br18_trueOut),
    .ins_valid (cond_br18_trueOut_valid),
    .ins_ready (cond_br18_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer44_outs),
    .outs_valid (buffer44_outs_valid),
    .outs_ready (buffer44_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer45(
    .ins (buffer44_outs),
    .ins_valid (buffer44_outs_valid),
    .ins_ready (buffer44_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer45_outs),
    .outs_valid (buffer45_outs_valid),
    .outs_ready (buffer45_outs_ready)
  );

  oehb_dataless buffer56(
    .ins_valid (cond_br24_trueOut_valid),
    .ins_ready (cond_br24_trueOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer56_outs_valid),
    .outs_ready (buffer56_outs_ready)
  );

  tehb_dataless buffer57(
    .ins_valid (buffer56_outs_valid),
    .ins_ready (buffer56_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer57_outs_valid),
    .outs_ready (buffer57_outs_ready)
  );

  source source2(
    .clk (clk),
    .rst (rst),
    .outs_valid (source2_outs_valid),
    .outs_ready (source2_outs_ready)
  );

  handshake_constant_3 #(.DATA_WIDTH(32)) constant6(
    .ctrl_valid (source2_outs_valid),
    .ctrl_ready (source2_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (constant6_outs),
    .outs_valid (constant6_outs_valid),
    .outs_ready (constant6_outs_ready)
  );

  trunci #(.INPUT_TYPE(32), .OUTPUT_TYPE(8)) trunci4(
    .ins (constant6_outs),
    .ins_valid (constant6_outs_valid),
    .ins_ready (constant6_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (trunci4_outs),
    .outs_valid (trunci4_outs_valid),
    .outs_ready (trunci4_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer62(
    .ins (cond_br20_falseOut),
    .ins_valid (cond_br20_falseOut_valid),
    .ins_ready (cond_br20_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer62_outs),
    .outs_valid (buffer62_outs_valid),
    .outs_ready (buffer62_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer63(
    .ins (buffer62_outs),
    .ins_valid (buffer62_outs_valid),
    .ins_ready (buffer62_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer63_outs),
    .outs_valid (buffer63_outs_valid),
    .outs_ready (buffer63_outs_ready)
  );

  addi #(.DATA_TYPE(8)) addi2(
    .lhs (buffer63_outs),
    .lhs_valid (buffer63_outs_valid),
    .lhs_ready (buffer63_outs_ready),
    .rhs (trunci4_outs),
    .rhs_valid (trunci4_outs_valid),
    .rhs_ready (trunci4_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (addi2_result),
    .result_valid (addi2_result_valid),
    .result_ready (addi2_result_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer60(
    .ins (cond_br25_falseOut),
    .ins_valid (cond_br25_falseOut_valid),
    .ins_ready (cond_br25_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer60_outs),
    .outs_valid (buffer60_outs_valid),
    .outs_ready (buffer60_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer61(
    .ins (buffer60_outs),
    .ins_valid (buffer60_outs_valid),
    .ins_ready (buffer60_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer61_outs),
    .outs_valid (buffer61_outs_valid),
    .outs_ready (buffer61_outs_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer66(
    .ins (cond_br22_falseOut),
    .ins_valid (cond_br22_falseOut_valid),
    .ins_ready (cond_br22_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer66_outs),
    .outs_valid (buffer66_outs_valid),
    .outs_ready (buffer66_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer67(
    .ins (buffer66_outs),
    .ins_valid (buffer66_outs_valid),
    .ins_ready (buffer66_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer67_outs),
    .outs_valid (buffer67_outs_valid),
    .outs_ready (buffer67_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer68(
    .ins (cond_br23_falseOut),
    .ins_valid (cond_br23_falseOut_valid),
    .ins_ready (cond_br23_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer68_outs),
    .outs_valid (buffer68_outs_valid),
    .outs_ready (buffer68_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer69(
    .ins (buffer68_outs),
    .ins_valid (buffer68_outs_valid),
    .ins_ready (buffer68_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer69_outs),
    .outs_valid (buffer69_outs_valid),
    .outs_ready (buffer69_outs_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer64(
    .ins (cond_br21_falseOut),
    .ins_valid (cond_br21_falseOut_valid),
    .ins_ready (cond_br21_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer64_outs),
    .outs_valid (buffer64_outs_valid),
    .outs_ready (buffer64_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer65(
    .ins (buffer64_outs),
    .ins_valid (buffer64_outs_valid),
    .ins_ready (buffer64_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer65_outs),
    .outs_valid (buffer65_outs_valid),
    .outs_ready (buffer65_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer58(
    .ins (cond_br18_falseOut),
    .ins_valid (cond_br18_falseOut_valid),
    .ins_ready (cond_br18_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer58_outs),
    .outs_valid (buffer58_outs_valid),
    .outs_ready (buffer58_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer59(
    .ins (buffer58_outs),
    .ins_valid (buffer58_outs_valid),
    .ins_ready (buffer58_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer59_outs),
    .outs_valid (buffer59_outs_valid),
    .outs_ready (buffer59_outs_ready)
  );

  oehb_dataless buffer70(
    .ins_valid (cond_br24_falseOut_valid),
    .ins_ready (cond_br24_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer70_outs_valid),
    .outs_ready (buffer70_outs_ready)
  );

  tehb_dataless buffer71(
    .ins_valid (buffer70_outs_valid),
    .ins_ready (buffer70_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs_valid (buffer71_outs_valid),
    .outs_ready (buffer71_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer72(
    .ins (cond_br3_falseOut),
    .ins_valid (cond_br3_falseOut_valid),
    .ins_ready (cond_br3_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer72_outs),
    .outs_valid (buffer72_outs_valid),
    .outs_ready (buffer72_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer73(
    .ins (buffer72_outs),
    .ins_valid (buffer72_outs_valid),
    .ins_ready (buffer72_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer73_outs),
    .outs_valid (buffer73_outs_valid),
    .outs_ready (buffer73_outs_ready)
  );

  oehb #(.DATA_TYPE(1)) buffer74(
    .ins (cond_br4_falseOut),
    .ins_valid (cond_br4_falseOut_valid),
    .ins_ready (cond_br4_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer74_outs),
    .outs_valid (buffer74_outs_valid),
    .outs_ready (buffer74_outs_ready)
  );

  tehb #(.DATA_TYPE(1)) buffer75(
    .ins (buffer74_outs),
    .ins_valid (buffer74_outs_valid),
    .ins_ready (buffer74_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer75_outs),
    .outs_valid (buffer75_outs_valid),
    .outs_ready (buffer75_outs_ready)
  );

  oehb #(.DATA_TYPE(8)) buffer76(
    .ins (cond_br5_falseOut),
    .ins_valid (cond_br5_falseOut_valid),
    .ins_ready (cond_br5_falseOut_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer76_outs),
    .outs_valid (buffer76_outs_valid),
    .outs_ready (buffer76_outs_ready)
  );

  tehb #(.DATA_TYPE(8)) buffer77(
    .ins (buffer76_outs),
    .ins_valid (buffer76_outs_valid),
    .ins_ready (buffer76_outs_ready),
    .clk (clk),
    .rst (rst),
    .outs (buffer77_outs),
    .outs_valid (buffer77_outs_valid),
    .outs_ready (buffer77_outs_ready)
  );

  selector #(.DATA_TYPE(8)) select1(
    .condition (buffer75_outs),
    .condition_valid (buffer75_outs_valid),
    .condition_ready (buffer75_outs_ready),
    .trueValue (buffer73_outs),
    .trueValue_valid (buffer73_outs_valid),
    .trueValue_ready (buffer73_outs_ready),
    .falseValue (buffer77_outs),
    .falseValue_valid (buffer77_outs_valid),
    .falseValue_ready (buffer77_outs_ready),
    .clk (clk),
    .rst (rst),
    .result (select1_result),
    .result_valid (select1_result_valid),
    .result_ready (select1_result_ready)
  );

endmodule
